module fsm1_route(
input GCLK_Pad,
input input1_Pad,
input input2_Pad,
input reset_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output output1_Pad);

wire net0_c1;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire reset_Pad;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire input1_Pad;
wire net58;
wire input2_Pad;
wire net59;
wire net60_c1;
wire output1_Pad;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire state_obs0_Pad;
wire net90_c1;
wire state_obs1_Pad;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire GCLK_Pad;
wire net207;

DFFT DFFT_61_state_obs0(net139,net80,net89_c1);
DFFT DFFT_56_state_obs1(net151,net88,net90_c1);
AND2T AND2T_9_n15(net102,net52,net76,net7_c1);
DFFT DFFT_51_output1(net101,net74,net60_c1);
NOTT NOTT_8_n14(net193,net45,net4_c1);
AND2T AND2T_11_n17(net203,net41,net79,net13_c1);
AND2T AND2T_21_n27(net115,net15,net54,net18_c1);
AND2T AND2T_13_n19(net100,net35,net23,net19_c1);
AND2T AND2T_30_n36(net147,net50,net87,net20_c1);
AND2T AND2T_15_n21(net163,net51,net83,net1_c1);
AND2T AND2T_24_n30(net148,net22,net75,net2_c1);
AND2T AND2T_16_n22(net167,net1,net49,net3_c1);
AND2T AND2T_18_n24(net127,net53,net63,net9_c1);
AND2T AND2T_19_n25(net99,net56,net43,net12_c1);
AND2T AND2T_28_n34(net194,net11,net85,net14_c1);
AND2T AND2T_29_n35(net199,net14,net8,net17_c1);
OR2T OR2T_20_n26(net116,net34,net33,net15_c1);
OR2T OR2T_22_n28(net125,net18,net12,net21_c1);
OR2T OR2T_23_n29(net126,net21,net64,net22_c1);
OR2T OR2T_26_n32(net187,net5,net78,net8_c1);
OR2T OR2T_27_n33(net200,net55,net25,net11_c1);
NOTT NOTT_10_n16(net191,net44,net10_c1);
NOTT NOTT_12_n18(net173,net40,net16_c1);
NOTT NOTT_14_n20(net98,net46,net0_c1);
NOTT NOTT_25_n31(net188,net38,net5_c1);
NOTT NOTT_17_n23(net164,net48,net6_c1);
DFFT DFFT_31__FBL_n124(net135,net2,net61_c1);
DFFT DFFT_32__FBL_n125(net205,net72,net62_c1);
DFFT DFFT_40__FPB_n133(net179,net66,net68_c1);
DFFT DFFT_41__FPB_n134(net177,net68,net71_c1);
DFFT DFFT_33__FPB_n126(net97,net17,net72_c1);
DFFT DFFT_50__FPB_n143(net111,net70,net74_c1);
DFFT DFFT_42__FPB_n135(net180,net71,net75_c1);
DFFT DFFT_34__FPB_n127(net136,net26,net76_c1);
DFFT DFFT_43__FPB_n136(net128,net31,net78_c1);
DFFT DFFT_35__FPB_n128(net206,net29,net79_c1);
DFFT DFFT_60__FPB_n153(net141,net77,net80_c1);
DFFT DFFT_52__FPB_n145(net204,net42,net81_c1);
DFFT DFFT_44__FPB_n137(net168,net27,net82_c1);
DFFT DFFT_36__FPB_n129(net96,net30,net83_c1);
DFFT DFFT_37__FPB_n130(net121,net28,net63_c1);
DFFT DFFT_53__FPB_n146(net192,net81,net84_c1);
DFFT DFFT_45__FPB_n138(net178,net82,net85_c1);
DFFT DFFT_38__FPB_n131(net95,net3,net64_c1);
DFFT DFFT_54__FPB_n147(net153,net84,net86_c1);
DFFT DFFT_46__FPB_n139(net154,net57,net87_c1);
DFFT DFFT_47__FPB_n140(net112,net37,net65_c1);
DFFT DFFT_39__FPB_n132(net174,net47,net66_c1);
DFFT DFFT_55__FPB_n148(net152,net86,net88_c1);
DFFT DFFT_48__FPB_n141(net94,net65,net67_c1);
DFFT DFFT_57__FPB_n150(net93,net20,net69_c1);
DFFT DFFT_49__FPB_n142(net122,net67,net70_c1);
DFFT DFFT_58__FPB_n151(net142,net69,net73_c1);
DFFT DFFT_59__FPB_n152(net140,net73,net77_c1);
SPLITT Split_62_n155(net58,net28_c1,net46_c1);
SPLITT Split_70_n163(net16,net27_c1,net47_c1);
SPLITT Split_63_n156(net59,net30_c1,net48_c1);
SPLITT Split_71_n164(net19,net31_c1,net49_c1);
SPLITT Split_64_n157(net4,net32_c1,net50_c1);
SPLITT Split_72_n165(net0,net33_c1,net51_c1);
SPLITT Split_65_n158(net32,net35_c1,net52_c1);
SPLITT Split_73_n166(net6,net34_c1,net53_c1);
SPLITT Split_66_n159(net7,net37_c1,net54_c1);
SPLITT Split_74_n167(net9,net36_c1,net55_c1);
SPLITT Split_67_n160(net10,net23_c1,net41_c1);
SPLITT Split_75_n168(net36,net38_c1,net56_c1);
SPLITT Split_68_n161(net13,net24_c1,net42_c1);
SPLITT Split_76_n169(net61,net39_c1,net57_c1);
SPLITT Split_69_n162(net24,net25_c1,net43_c1);
SPLITT Split_77_n170(net39,net26_c1,net44_c1);
SPLITT Split_78_n171(net62,net29_c1,net45_c1);
SPLITT SplitCLK_4_55(net201,net206_c1,net205_c1);
SPLITT SplitCLK_0_56(net202,net203_c1,net204_c1);
SPLITT SplitCLK_0_57(net195,net202_c1,net201_c1);
SPLITT SplitCLK_4_58(net198,net199_c1,net200_c1);
SPLITT SplitCLK_4_59(net196,net197_c1,net198_c1);
SPLITT SplitCLK_4_60(net181,net195_c1,net196_c1);
SPLITT SplitCLK_4_61(net189,net193_c1,net194_c1);
SPLITT SplitCLK_4_62(net190,net192_c1,net191_c1);
SPLITT SplitCLK_6_63(net183,net189_c1,net190_c1);
SPLITT SplitCLK_4_64(net186,net188_c1,net187_c1);
SPLITT SplitCLK_4_65(net184,net185_c1,net186_c1);
SPLITT SplitCLK_6_66(net182,net184_c1,net183_c1);
SPLITT SplitCLK_6_67(net155,net181_c1,net182_c1);
SPLITT SplitCLK_4_68(net175,net179_c1,net180_c1);
SPLITT SplitCLK_4_69(net176,net178_c1,net177_c1);
SPLITT SplitCLK_6_70(net169,net175_c1,net176_c1);
SPLITT SplitCLK_4_71(net172,net174_c1,net173_c1);
SPLITT SplitCLK_2_72(net170,net171_c1,net172_c1);
SPLITT SplitCLK_0_73(net157,net169_c1,net170_c1);
SPLITT SplitCLK_4_74(net166,net167_c1,net168_c1);
SPLITT SplitCLK_0_75(net159,net165_c1,net166_c1);
SPLITT SplitCLK_4_76(net162,net163_c1,net164_c1);
SPLITT SplitCLK_4_77(net160,net161_c1,net162_c1);
SPLITT SplitCLK_2_78(net158,net160_c1,net159_c1);
SPLITT SplitCLK_4_79(net156,net158_c1,net157_c1);
SPLITT SplitCLK_0_80(net91,net155_c1,net156_c1);
SPLITT SplitCLK_4_81(net149,net153_c1,net154_c1);
SPLITT SplitCLK_0_82(net150,net151_c1,net152_c1);
SPLITT SplitCLK_0_83(net143,net150_c1,net149_c1);
SPLITT SplitCLK_4_84(net146,net148_c1,net147_c1);
SPLITT SplitCLK_4_85(net144,net145_c1,net146_c1);
SPLITT SplitCLK_0_86(net129,net143_c1,net144_c1);
SPLITT SplitCLK_4_87(net137,net141_c1,net142_c1);
SPLITT SplitCLK_4_88(net138,net139_c1,net140_c1);
SPLITT SplitCLK_6_89(net131,net137_c1,net138_c1);
SPLITT SplitCLK_4_90(net134,net135_c1,net136_c1);
SPLITT SplitCLK_4_91(net132,net133_c1,net134_c1);
SPLITT SplitCLK_2_92(net130,net132_c1,net131_c1);
SPLITT SplitCLK_6_93(net103,net129_c1,net130_c1);
SPLITT SplitCLK_4_94(net123,net128_c1,net127_c1);
SPLITT SplitCLK_4_95(net124,net125_c1,net126_c1);
SPLITT SplitCLK_4_96(net117,net124_c1,net123_c1);
SPLITT SplitCLK_4_97(net120,net121_c1,net122_c1);
SPLITT SplitCLK_4_98(net118,net119_c1,net120_c1);
SPLITT SplitCLK_0_99(net105,net117_c1,net118_c1);
SPLITT SplitCLK_4_100(net114,net115_c1,net116_c1);
SPLITT SplitCLK_6_101(net107,net114_c1,net113_c1);
SPLITT SplitCLK_4_102(net110,net112_c1,net111_c1);
SPLITT SplitCLK_2_103(net108,net109_c1,net110_c1);
SPLITT SplitCLK_4_104(net106,net107_c1,net108_c1);
SPLITT SplitCLK_4_105(net104,net106_c1,net105_c1);
SPLITT SplitCLK_2_106(net92,net104_c1,net103_c1);
wire dummy0;
SPLITT SplitCLK_2_107(net133,net102_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_2_108(net109,net101_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_109(net185,net100_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_110(net113,net99_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_111(net161,net98_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_2_112(net197,net97_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_2_113(net171,net96_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_2_114(net165,net95_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_2_115(net119,net94_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_2_116(net145,net93_c1,dummy9);
SPLITT SplitCLK_0_117(net207,net91_c1,net92_c1);
INTERCONNECT NOTT_14_n20_Split_72_n165(net0_c1,net0);
INTERCONNECT AND2T_15_n21_AND2T_16_n22(net1_c1,net1);
INTERCONNECT AND2T_24_n30_DFFT_31__FBL_n124(net2_c1,net2);
INTERCONNECT AND2T_16_n22_DFFT_38__FPB_n131(net3_c1,net3);
INTERCONNECT NOTT_8_n14_Split_64_n157(net4_c1,net4);
INTERCONNECT NOTT_25_n31_OR2T_26_n32(net5_c1,net5);
INTERCONNECT NOTT_17_n23_Split_73_n166(net6_c1,net6);
INTERCONNECT AND2T_9_n15_Split_66_n159(net7_c1,net7);
INTERCONNECT OR2T_26_n32_AND2T_29_n35(net8_c1,net8);
INTERCONNECT AND2T_18_n24_Split_74_n167(net9_c1,net9);
INTERCONNECT NOTT_10_n16_Split_67_n160(net10_c1,net10);
INTERCONNECT OR2T_27_n33_AND2T_28_n34(net11_c1,net11);
INTERCONNECT AND2T_19_n25_OR2T_22_n28(net12_c1,net12);
INTERCONNECT AND2T_11_n17_Split_68_n161(net13_c1,net13);
INTERCONNECT AND2T_28_n34_AND2T_29_n35(net14_c1,net14);
INTERCONNECT OR2T_20_n26_AND2T_21_n27(net15_c1,net15);
INTERCONNECT NOTT_12_n18_Split_70_n163(net16_c1,net16);
INTERCONNECT AND2T_29_n35_DFFT_33__FPB_n126(net17_c1,net17);
INTERCONNECT AND2T_21_n27_OR2T_22_n28(net18_c1,net18);
INTERCONNECT AND2T_13_n19_Split_71_n164(net19_c1,net19);
INTERCONNECT AND2T_30_n36_DFFT_57__FPB_n150(net20_c1,net20);
INTERCONNECT OR2T_22_n28_OR2T_23_n29(net21_c1,net21);
INTERCONNECT OR2T_23_n29_AND2T_24_n30(net22_c1,net22);
INTERCONNECT Split_67_n160_AND2T_13_n19(net23_c1,net23);
INTERCONNECT Split_68_n161_Split_69_n162(net24_c1,net24);
INTERCONNECT Split_69_n162_OR2T_27_n33(net25_c1,net25);
INTERCONNECT Split_77_n170_DFFT_34__FPB_n127(net26_c1,net26);
INTERCONNECT Split_70_n163_DFFT_44__FPB_n137(net27_c1,net27);
INTERCONNECT Split_62_n155_DFFT_37__FPB_n130(net28_c1,net28);
INTERCONNECT Split_78_n171_DFFT_35__FPB_n128(net29_c1,net29);
INTERCONNECT Split_63_n156_DFFT_36__FPB_n129(net30_c1,net30);
INTERCONNECT Split_71_n164_DFFT_43__FPB_n136(net31_c1,net31);
INTERCONNECT Split_64_n157_Split_65_n158(net32_c1,net32);
INTERCONNECT Split_72_n165_OR2T_20_n26(net33_c1,net33);
INTERCONNECT Split_73_n166_OR2T_20_n26(net34_c1,net34);
INTERCONNECT Split_65_n158_AND2T_13_n19(net35_c1,net35);
INTERCONNECT Split_74_n167_Split_75_n168(net36_c1,net36);
INTERCONNECT Split_66_n159_DFFT_47__FPB_n140(net37_c1,net37);
INTERCONNECT Split_75_n168_NOTT_25_n31(net38_c1,net38);
INTERCONNECT Split_76_n169_Split_77_n170(net39_c1,net39);
INTERCONNECT reset_Pad_NOTT_12_n18(reset_Pad,net40);
INTERCONNECT Split_67_n160_AND2T_11_n17(net41_c1,net41);
INTERCONNECT Split_68_n161_DFFT_52__FPB_n145(net42_c1,net42);
INTERCONNECT Split_69_n162_AND2T_19_n25(net43_c1,net43);
INTERCONNECT Split_77_n170_NOTT_10_n16(net44_c1,net44);
INTERCONNECT Split_78_n171_NOTT_8_n14(net45_c1,net45);
INTERCONNECT Split_62_n155_NOTT_14_n20(net46_c1,net46);
INTERCONNECT Split_70_n163_DFFT_39__FPB_n132(net47_c1,net47);
INTERCONNECT Split_63_n156_NOTT_17_n23(net48_c1,net48);
INTERCONNECT Split_71_n164_AND2T_16_n22(net49_c1,net49);
INTERCONNECT Split_64_n157_AND2T_30_n36(net50_c1,net50);
INTERCONNECT Split_72_n165_AND2T_15_n21(net51_c1,net51);
INTERCONNECT Split_65_n158_AND2T_9_n15(net52_c1,net52);
INTERCONNECT Split_73_n166_AND2T_18_n24(net53_c1,net53);
INTERCONNECT Split_66_n159_AND2T_21_n27(net54_c1,net54);
INTERCONNECT Split_74_n167_OR2T_27_n33(net55_c1,net55);
INTERCONNECT Split_75_n168_AND2T_19_n25(net56_c1,net56);
INTERCONNECT Split_76_n169_DFFT_46__FPB_n139(net57_c1,net57);
INTERCONNECT input1_Pad_Split_62_n155(input1_Pad,net58);
INTERCONNECT input2_Pad_Split_63_n156(input2_Pad,net59);
INTERCONNECT DFFT_51_output1_output1_Pad(net60_c1,output1_Pad);
INTERCONNECT DFFT_31__FBL_n124_Split_76_n169(net61_c1,net61);
INTERCONNECT DFFT_32__FBL_n125_Split_78_n171(net62_c1,net62);
INTERCONNECT DFFT_37__FPB_n130_AND2T_18_n24(net63_c1,net63);
INTERCONNECT DFFT_38__FPB_n131_OR2T_23_n29(net64_c1,net64);
INTERCONNECT DFFT_47__FPB_n140_DFFT_48__FPB_n141(net65_c1,net65);
INTERCONNECT DFFT_39__FPB_n132_DFFT_40__FPB_n133(net66_c1,net66);
INTERCONNECT DFFT_48__FPB_n141_DFFT_49__FPB_n142(net67_c1,net67);
INTERCONNECT DFFT_40__FPB_n133_DFFT_41__FPB_n134(net68_c1,net68);
INTERCONNECT DFFT_57__FPB_n150_DFFT_58__FPB_n151(net69_c1,net69);
INTERCONNECT DFFT_49__FPB_n142_DFFT_50__FPB_n143(net70_c1,net70);
INTERCONNECT DFFT_41__FPB_n134_DFFT_42__FPB_n135(net71_c1,net71);
INTERCONNECT DFFT_33__FPB_n126_DFFT_32__FBL_n125(net72_c1,net72);
INTERCONNECT DFFT_58__FPB_n151_DFFT_59__FPB_n152(net73_c1,net73);
INTERCONNECT DFFT_50__FPB_n143_DFFT_51_output1(net74_c1,net74);
INTERCONNECT DFFT_42__FPB_n135_AND2T_24_n30(net75_c1,net75);
INTERCONNECT DFFT_34__FPB_n127_AND2T_9_n15(net76_c1,net76);
INTERCONNECT DFFT_59__FPB_n152_DFFT_60__FPB_n153(net77_c1,net77);
INTERCONNECT DFFT_43__FPB_n136_OR2T_26_n32(net78_c1,net78);
INTERCONNECT DFFT_35__FPB_n128_AND2T_11_n17(net79_c1,net79);
INTERCONNECT DFFT_60__FPB_n153_DFFT_61_state_obs0(net80_c1,net80);
INTERCONNECT DFFT_52__FPB_n145_DFFT_53__FPB_n146(net81_c1,net81);
INTERCONNECT DFFT_44__FPB_n137_DFFT_45__FPB_n138(net82_c1,net82);
INTERCONNECT DFFT_36__FPB_n129_AND2T_15_n21(net83_c1,net83);
INTERCONNECT DFFT_53__FPB_n146_DFFT_54__FPB_n147(net84_c1,net84);
INTERCONNECT DFFT_45__FPB_n138_AND2T_28_n34(net85_c1,net85);
INTERCONNECT DFFT_54__FPB_n147_DFFT_55__FPB_n148(net86_c1,net86);
INTERCONNECT DFFT_46__FPB_n139_AND2T_30_n36(net87_c1,net87);
INTERCONNECT DFFT_55__FPB_n148_DFFT_56_state_obs1(net88_c1,net88);
INTERCONNECT DFFT_61_state_obs0_state_obs0_Pad(net89_c1,state_obs0_Pad);
INTERCONNECT DFFT_56_state_obs1_state_obs1_Pad(net90_c1,state_obs1_Pad);
INTERCONNECT SplitCLK_0_117_SplitCLK_0_80(net91_c1,net91);
INTERCONNECT SplitCLK_0_117_SplitCLK_2_106(net92_c1,net92);
INTERCONNECT SplitCLK_2_116_DFFT_57__FPB_n150(net93_c1,net93);
INTERCONNECT SplitCLK_2_115_DFFT_48__FPB_n141(net94_c1,net94);
INTERCONNECT SplitCLK_2_114_DFFT_38__FPB_n131(net95_c1,net95);
INTERCONNECT SplitCLK_2_113_DFFT_36__FPB_n129(net96_c1,net96);
INTERCONNECT SplitCLK_2_112_DFFT_33__FPB_n126(net97_c1,net97);
INTERCONNECT SplitCLK_2_111_NOTT_14_n20(net98_c1,net98);
INTERCONNECT SplitCLK_2_110_AND2T_19_n25(net99_c1,net99);
INTERCONNECT SplitCLK_2_109_AND2T_13_n19(net100_c1,net100);
INTERCONNECT SplitCLK_2_108_DFFT_51_output1(net101_c1,net101);
INTERCONNECT SplitCLK_2_107_AND2T_9_n15(net102_c1,net102);
INTERCONNECT SplitCLK_2_106_SplitCLK_6_93(net103_c1,net103);
INTERCONNECT SplitCLK_2_106_SplitCLK_4_105(net104_c1,net104);
INTERCONNECT SplitCLK_4_105_SplitCLK_0_99(net105_c1,net105);
INTERCONNECT SplitCLK_4_105_SplitCLK_4_104(net106_c1,net106);
INTERCONNECT SplitCLK_4_104_SplitCLK_6_101(net107_c1,net107);
INTERCONNECT SplitCLK_4_104_SplitCLK_2_103(net108_c1,net108);
INTERCONNECT SplitCLK_2_103_SplitCLK_2_108(net109_c1,net109);
INTERCONNECT SplitCLK_2_103_SplitCLK_4_102(net110_c1,net110);
INTERCONNECT SplitCLK_4_102_DFFT_50__FPB_n143(net111_c1,net111);
INTERCONNECT SplitCLK_4_102_DFFT_47__FPB_n140(net112_c1,net112);
INTERCONNECT SplitCLK_6_101_SplitCLK_2_110(net113_c1,net113);
INTERCONNECT SplitCLK_6_101_SplitCLK_4_100(net114_c1,net114);
INTERCONNECT SplitCLK_4_100_AND2T_21_n27(net115_c1,net115);
INTERCONNECT SplitCLK_4_100_OR2T_20_n26(net116_c1,net116);
INTERCONNECT SplitCLK_0_99_SplitCLK_4_96(net117_c1,net117);
INTERCONNECT SplitCLK_0_99_SplitCLK_4_98(net118_c1,net118);
INTERCONNECT SplitCLK_4_98_SplitCLK_2_115(net119_c1,net119);
INTERCONNECT SplitCLK_4_98_SplitCLK_4_97(net120_c1,net120);
INTERCONNECT SplitCLK_4_97_DFFT_37__FPB_n130(net121_c1,net121);
INTERCONNECT SplitCLK_4_97_DFFT_49__FPB_n142(net122_c1,net122);
INTERCONNECT SplitCLK_4_96_SplitCLK_4_94(net123_c1,net123);
INTERCONNECT SplitCLK_4_96_SplitCLK_4_95(net124_c1,net124);
INTERCONNECT SplitCLK_4_95_OR2T_22_n28(net125_c1,net125);
INTERCONNECT SplitCLK_4_95_OR2T_23_n29(net126_c1,net126);
INTERCONNECT SplitCLK_4_94_AND2T_18_n24(net127_c1,net127);
INTERCONNECT SplitCLK_4_94_DFFT_43__FPB_n136(net128_c1,net128);
INTERCONNECT SplitCLK_6_93_SplitCLK_0_86(net129_c1,net129);
INTERCONNECT SplitCLK_6_93_SplitCLK_2_92(net130_c1,net130);
INTERCONNECT SplitCLK_2_92_SplitCLK_6_89(net131_c1,net131);
INTERCONNECT SplitCLK_2_92_SplitCLK_4_91(net132_c1,net132);
INTERCONNECT SplitCLK_4_91_SplitCLK_2_107(net133_c1,net133);
INTERCONNECT SplitCLK_4_91_SplitCLK_4_90(net134_c1,net134);
INTERCONNECT SplitCLK_4_90_DFFT_31__FBL_n124(net135_c1,net135);
INTERCONNECT SplitCLK_4_90_DFFT_34__FPB_n127(net136_c1,net136);
INTERCONNECT SplitCLK_6_89_SplitCLK_4_87(net137_c1,net137);
INTERCONNECT SplitCLK_6_89_SplitCLK_4_88(net138_c1,net138);
INTERCONNECT SplitCLK_4_88_DFFT_61_state_obs0(net139_c1,net139);
INTERCONNECT SplitCLK_4_88_DFFT_59__FPB_n152(net140_c1,net140);
INTERCONNECT SplitCLK_4_87_DFFT_60__FPB_n153(net141_c1,net141);
INTERCONNECT SplitCLK_4_87_DFFT_58__FPB_n151(net142_c1,net142);
INTERCONNECT SplitCLK_0_86_SplitCLK_0_83(net143_c1,net143);
INTERCONNECT SplitCLK_0_86_SplitCLK_4_85(net144_c1,net144);
INTERCONNECT SplitCLK_4_85_SplitCLK_2_116(net145_c1,net145);
INTERCONNECT SplitCLK_4_85_SplitCLK_4_84(net146_c1,net146);
INTERCONNECT SplitCLK_4_84_AND2T_30_n36(net147_c1,net147);
INTERCONNECT SplitCLK_4_84_AND2T_24_n30(net148_c1,net148);
INTERCONNECT SplitCLK_0_83_SplitCLK_4_81(net149_c1,net149);
INTERCONNECT SplitCLK_0_83_SplitCLK_0_82(net150_c1,net150);
INTERCONNECT SplitCLK_0_82_DFFT_56_state_obs1(net151_c1,net151);
INTERCONNECT SplitCLK_0_82_DFFT_55__FPB_n148(net152_c1,net152);
INTERCONNECT SplitCLK_4_81_DFFT_54__FPB_n147(net153_c1,net153);
INTERCONNECT SplitCLK_4_81_DFFT_46__FPB_n139(net154_c1,net154);
INTERCONNECT SplitCLK_0_80_SplitCLK_6_67(net155_c1,net155);
INTERCONNECT SplitCLK_0_80_SplitCLK_4_79(net156_c1,net156);
INTERCONNECT SplitCLK_4_79_SplitCLK_0_73(net157_c1,net157);
INTERCONNECT SplitCLK_4_79_SplitCLK_2_78(net158_c1,net158);
INTERCONNECT SplitCLK_2_78_SplitCLK_0_75(net159_c1,net159);
INTERCONNECT SplitCLK_2_78_SplitCLK_4_77(net160_c1,net160);
INTERCONNECT SplitCLK_4_77_SplitCLK_2_111(net161_c1,net161);
INTERCONNECT SplitCLK_4_77_SplitCLK_4_76(net162_c1,net162);
INTERCONNECT SplitCLK_4_76_AND2T_15_n21(net163_c1,net163);
INTERCONNECT SplitCLK_4_76_NOTT_17_n23(net164_c1,net164);
INTERCONNECT SplitCLK_0_75_SplitCLK_2_114(net165_c1,net165);
INTERCONNECT SplitCLK_0_75_SplitCLK_4_74(net166_c1,net166);
INTERCONNECT SplitCLK_4_74_AND2T_16_n22(net167_c1,net167);
INTERCONNECT SplitCLK_4_74_DFFT_44__FPB_n137(net168_c1,net168);
INTERCONNECT SplitCLK_0_73_SplitCLK_6_70(net169_c1,net169);
INTERCONNECT SplitCLK_0_73_SplitCLK_2_72(net170_c1,net170);
INTERCONNECT SplitCLK_2_72_SplitCLK_2_113(net171_c1,net171);
INTERCONNECT SplitCLK_2_72_SplitCLK_4_71(net172_c1,net172);
INTERCONNECT SplitCLK_4_71_NOTT_12_n18(net173_c1,net173);
INTERCONNECT SplitCLK_4_71_DFFT_39__FPB_n132(net174_c1,net174);
INTERCONNECT SplitCLK_6_70_SplitCLK_4_68(net175_c1,net175);
INTERCONNECT SplitCLK_6_70_SplitCLK_4_69(net176_c1,net176);
INTERCONNECT SplitCLK_4_69_DFFT_41__FPB_n134(net177_c1,net177);
INTERCONNECT SplitCLK_4_69_DFFT_45__FPB_n138(net178_c1,net178);
INTERCONNECT SplitCLK_4_68_DFFT_40__FPB_n133(net179_c1,net179);
INTERCONNECT SplitCLK_4_68_DFFT_42__FPB_n135(net180_c1,net180);
INTERCONNECT SplitCLK_6_67_SplitCLK_4_60(net181_c1,net181);
INTERCONNECT SplitCLK_6_67_SplitCLK_6_66(net182_c1,net182);
INTERCONNECT SplitCLK_6_66_SplitCLK_6_63(net183_c1,net183);
INTERCONNECT SplitCLK_6_66_SplitCLK_4_65(net184_c1,net184);
INTERCONNECT SplitCLK_4_65_SplitCLK_2_109(net185_c1,net185);
INTERCONNECT SplitCLK_4_65_SplitCLK_4_64(net186_c1,net186);
INTERCONNECT SplitCLK_4_64_OR2T_26_n32(net187_c1,net187);
INTERCONNECT SplitCLK_4_64_NOTT_25_n31(net188_c1,net188);
INTERCONNECT SplitCLK_6_63_SplitCLK_4_61(net189_c1,net189);
INTERCONNECT SplitCLK_6_63_SplitCLK_4_62(net190_c1,net190);
INTERCONNECT SplitCLK_4_62_NOTT_10_n16(net191_c1,net191);
INTERCONNECT SplitCLK_4_62_DFFT_53__FPB_n146(net192_c1,net192);
INTERCONNECT SplitCLK_4_61_NOTT_8_n14(net193_c1,net193);
INTERCONNECT SplitCLK_4_61_AND2T_28_n34(net194_c1,net194);
INTERCONNECT SplitCLK_4_60_SplitCLK_0_57(net195_c1,net195);
INTERCONNECT SplitCLK_4_60_SplitCLK_4_59(net196_c1,net196);
INTERCONNECT SplitCLK_4_59_SplitCLK_2_112(net197_c1,net197);
INTERCONNECT SplitCLK_4_59_SplitCLK_4_58(net198_c1,net198);
INTERCONNECT SplitCLK_4_58_AND2T_29_n35(net199_c1,net199);
INTERCONNECT SplitCLK_4_58_OR2T_27_n33(net200_c1,net200);
INTERCONNECT SplitCLK_0_57_SplitCLK_4_55(net201_c1,net201);
INTERCONNECT SplitCLK_0_57_SplitCLK_0_56(net202_c1,net202);
INTERCONNECT SplitCLK_0_56_AND2T_11_n17(net203_c1,net203);
INTERCONNECT SplitCLK_0_56_DFFT_52__FPB_n145(net204_c1,net204);
INTERCONNECT SplitCLK_4_55_DFFT_32__FBL_n125(net205_c1,net205);
INTERCONNECT SplitCLK_4_55_DFFT_35__FPB_n128(net206_c1,net206);
INTERCONNECT GCLK_Pad_SplitCLK_0_117(GCLK_Pad,net207);

endmodule
