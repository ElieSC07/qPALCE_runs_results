module ID4s_route(
input GCLK_Pad,
input D0_Pad,
input D1_Pad,
input D2_Pad,
input D3_Pad,
input X0_Pad,
input X1_Pad,
input X2_Pad,
input X3_Pad,
output Q0_Pad,
output Q1_Pad,
output R0_Pad,
output Q2_Pad,
output R1_Pad,
output Q3_Pad,
output R2_Pad,
output R3_Pad);

wire D0_Pad;
wire net0;
wire D1_Pad;
wire net1;
wire D2_Pad;
wire net2;
wire D3_Pad;
wire net3;
wire net4_c1;
wire Q0_Pad;
wire net5_c1;
wire Q1_Pad;
wire net6_c1;
wire R0_Pad;
wire net7_c1;
wire Q2_Pad;
wire net8_c1;
wire R1_Pad;
wire net9_c1;
wire Q3_Pad;
wire net10_c1;
wire R2_Pad;
wire net11_c1;
wire R3_Pad;
wire X0_Pad;
wire net12;
wire X1_Pad;
wire net13;
wire X2_Pad;
wire net14;
wire X3_Pad;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire net486_c1;
wire net486;
wire net487_c1;
wire net487;
wire net488_c1;
wire net488;
wire net489_c1;
wire net489;
wire net490_c1;
wire net490;
wire net491_c1;
wire net491;
wire net492_c1;
wire net492;
wire net493_c1;
wire net493;
wire net494_c1;
wire net494;
wire net495_c1;
wire net495;
wire net496_c1;
wire net496;
wire net497_c1;
wire net497;
wire net498_c1;
wire net498;
wire net499_c1;
wire net499;
wire net500_c1;
wire net500;
wire net501_c1;
wire net501;
wire net502_c1;
wire net502;
wire net503_c1;
wire net503;
wire net504_c1;
wire net504;
wire net505_c1;
wire net505;
wire net506_c1;
wire net506;
wire net507_c1;
wire net507;
wire net508_c1;
wire net508;
wire net509_c1;
wire net509;
wire net510_c1;
wire net510;
wire net511_c1;
wire net511;
wire net512_c1;
wire net512;
wire net513_c1;
wire net513;
wire net514_c1;
wire net514;
wire net515_c1;
wire net515;
wire net516_c1;
wire net516;
wire net517_c1;
wire net517;
wire net518_c1;
wire net518;
wire net519_c1;
wire net519;
wire net520_c1;
wire net520;
wire net521_c1;
wire net521;
wire net522_c1;
wire net522;
wire net523_c1;
wire net523;
wire net524_c1;
wire net524;
wire net525_c1;
wire net525;
wire net526_c1;
wire net526;
wire net527_c1;
wire net527;
wire net528_c1;
wire net528;
wire net529_c1;
wire net529;
wire net530_c1;
wire net530;
wire net531_c1;
wire net531;
wire net532_c1;
wire net532;
wire net533_c1;
wire net533;
wire net534_c1;
wire net534;
wire net535_c1;
wire net535;
wire net536_c1;
wire net536;
wire net537_c1;
wire net537;
wire net538_c1;
wire net538;
wire net539_c1;
wire net539;
wire net540_c1;
wire net540;
wire net541_c1;
wire net541;
wire net542_c1;
wire net542;
wire net543_c1;
wire net543;
wire net544_c1;
wire net544;
wire net545_c1;
wire net545;
wire net546_c1;
wire net546;
wire net547_c1;
wire net547;
wire net548_c1;
wire net548;
wire net549_c1;
wire net549;
wire net550_c1;
wire net550;
wire net551_c1;
wire net551;
wire net552_c1;
wire net552;
wire net553_c1;
wire net553;
wire net554_c1;
wire net554;
wire net555_c1;
wire net555;
wire net556_c1;
wire net556;
wire net557_c1;
wire net557;
wire net558_c1;
wire net558;
wire net559_c1;
wire net559;
wire net560_c1;
wire net560;
wire net561_c1;
wire net561;
wire net562_c1;
wire net562;
wire net563_c1;
wire net563;
wire net564_c1;
wire net564;
wire net565_c1;
wire net565;
wire net566_c1;
wire net566;
wire net567_c1;
wire net567;
wire net568_c1;
wire net568;
wire net569_c1;
wire net569;
wire net570_c1;
wire net570;
wire net571_c1;
wire net571;
wire net572_c1;
wire net572;
wire net573_c1;
wire net573;
wire net574_c1;
wire net574;
wire net575_c1;
wire net575;
wire net576_c1;
wire net576;
wire net577_c1;
wire net577;
wire net578_c1;
wire net578;
wire net579_c1;
wire net579;
wire net580_c1;
wire net580;
wire net581_c1;
wire net581;
wire net582_c1;
wire net582;
wire net583_c1;
wire net583;
wire net584_c1;
wire net584;
wire net585_c1;
wire net585;
wire net586_c1;
wire net586;
wire net587_c1;
wire net587;
wire net588_c1;
wire net588;
wire net589_c1;
wire net589;
wire net590_c1;
wire net590;
wire net591_c1;
wire net591;
wire net592_c1;
wire net592;
wire net593_c1;
wire net593;
wire net594_c1;
wire net594;
wire net595_c1;
wire net595;
wire net596_c1;
wire net596;
wire net597_c1;
wire net597;
wire net598_c1;
wire net598;
wire net599_c1;
wire net599;
wire net600_c1;
wire net600;
wire net601_c1;
wire net601;
wire net602_c1;
wire net602;
wire net603_c1;
wire net603;
wire net604_c1;
wire net604;
wire net605_c1;
wire net605;
wire net606_c1;
wire net606;
wire net607_c1;
wire net607;
wire net608_c1;
wire net608;
wire net609_c1;
wire net609;
wire net610_c1;
wire net610;
wire net611_c1;
wire net611;
wire net612_c1;
wire net612;
wire net613_c1;
wire net613;
wire net614_c1;
wire net614;
wire net615_c1;
wire net615;
wire net616_c1;
wire net616;
wire net617_c1;
wire net617;
wire net618_c1;
wire net618;
wire net619_c1;
wire net619;
wire net620_c1;
wire net620;
wire net621_c1;
wire net621;
wire net622_c1;
wire net622;
wire net623_c1;
wire net623;
wire net624_c1;
wire net624;
wire net625_c1;
wire net625;
wire net626_c1;
wire net626;
wire net627_c1;
wire net627;
wire net628_c1;
wire net628;
wire net629_c1;
wire net629;
wire net630_c1;
wire net630;
wire net631_c1;
wire net631;
wire net632_c1;
wire net632;
wire net633_c1;
wire net633;
wire net634_c1;
wire net634;
wire net635_c1;
wire net635;
wire net636_c1;
wire net636;
wire net637_c1;
wire net637;
wire net638_c1;
wire net638;
wire net639_c1;
wire net639;
wire net640_c1;
wire net640;
wire net641_c1;
wire net641;
wire net642_c1;
wire net642;
wire net643_c1;
wire net643;
wire net644_c1;
wire net644;
wire net645_c1;
wire net645;
wire net646_c1;
wire net646;
wire net647_c1;
wire net647;
wire net648_c1;
wire net648;
wire net649_c1;
wire net649;
wire net650_c1;
wire net650;
wire net651_c1;
wire net651;
wire net652_c1;
wire net652;
wire net653_c1;
wire net653;
wire net654_c1;
wire net654;
wire net655_c1;
wire net655;
wire net656_c1;
wire net656;
wire net657_c1;
wire net657;
wire net658_c1;
wire net658;
wire net659_c1;
wire net659;
wire net660_c1;
wire net660;
wire net661_c1;
wire net661;
wire net662_c1;
wire net662;
wire net663_c1;
wire net663;
wire net664_c1;
wire net664;
wire net665_c1;
wire net665;
wire net666_c1;
wire net666;
wire net667_c1;
wire net667;
wire net668_c1;
wire net668;
wire net669_c1;
wire net669;
wire net670_c1;
wire net670;
wire net671_c1;
wire net671;
wire net672_c1;
wire net672;
wire net673_c1;
wire net673;
wire net674_c1;
wire net674;
wire net675_c1;
wire net675;
wire net676_c1;
wire net676;
wire net677_c1;
wire net677;
wire net678_c1;
wire net678;
wire net679_c1;
wire net679;
wire net680_c1;
wire net680;
wire net681_c1;
wire net681;
wire net682_c1;
wire net682;
wire net683_c1;
wire net683;
wire net684_c1;
wire net684;
wire net685_c1;
wire net685;
wire net686_c1;
wire net686;
wire net687_c1;
wire net687;
wire net688_c1;
wire net688;
wire net689_c1;
wire net689;
wire net690_c1;
wire net690;
wire net691_c1;
wire net691;
wire net692_c1;
wire net692;
wire net693_c1;
wire net693;
wire net694_c1;
wire net694;
wire net695_c1;
wire net695;
wire net696_c1;
wire net696;
wire net697_c1;
wire net697;
wire net698_c1;
wire net698;
wire net699_c1;
wire net699;
wire net700_c1;
wire net700;
wire net701_c1;
wire net701;
wire net702_c1;
wire net702;
wire net703_c1;
wire net703;
wire net704_c1;
wire net704;
wire net705_c1;
wire net705;
wire net706_c1;
wire net706;
wire net707_c1;
wire net707;
wire net708_c1;
wire net708;
wire net709_c1;
wire net709;
wire net710_c1;
wire net710;
wire net711_c1;
wire net711;
wire net712_c1;
wire net712;
wire net713_c1;
wire net713;
wire net714_c1;
wire net714;
wire net715_c1;
wire net715;
wire net716_c1;
wire net716;
wire net717_c1;
wire net717;
wire net718_c1;
wire net718;
wire net719_c1;
wire net719;
wire net720_c1;
wire net720;
wire net721_c1;
wire net721;
wire net722_c1;
wire net722;
wire net723_c1;
wire net723;
wire net724_c1;
wire net724;
wire net725_c1;
wire net725;
wire net726_c1;
wire net726;
wire net727_c1;
wire net727;
wire net728_c1;
wire net728;
wire net729_c1;
wire net729;
wire net730_c1;
wire net730;
wire net731_c1;
wire net731;
wire net732_c1;
wire net732;
wire net733_c1;
wire net733;
wire net734_c1;
wire net734;
wire net735_c1;
wire net735;
wire net736_c1;
wire net736;
wire net737_c1;
wire net737;
wire net738_c1;
wire net738;
wire net739_c1;
wire net739;
wire net740_c1;
wire net740;
wire net741_c1;
wire net741;
wire net742_c1;
wire net742;
wire net743_c1;
wire net743;
wire net744_c1;
wire net744;
wire net745_c1;
wire net745;
wire net746_c1;
wire net746;
wire net747_c1;
wire net747;
wire net748_c1;
wire net748;
wire net749_c1;
wire net749;
wire net750_c1;
wire net750;
wire net751_c1;
wire net751;
wire net752_c1;
wire net752;
wire net753_c1;
wire net753;
wire net754_c1;
wire net754;
wire net755_c1;
wire net755;
wire net756_c1;
wire net756;
wire net757_c1;
wire net757;
wire net758_c1;
wire net758;
wire net759_c1;
wire net759;
wire net760_c1;
wire net760;
wire net761_c1;
wire net761;
wire net762_c1;
wire net762;
wire net763_c1;
wire net763;
wire net764_c1;
wire net764;
wire net765_c1;
wire net765;
wire net766_c1;
wire net766;
wire net767_c1;
wire net767;
wire net768_c1;
wire net768;
wire net769_c1;
wire net769;
wire net770_c1;
wire net770;
wire net771_c1;
wire net771;
wire net772_c1;
wire net772;
wire net773_c1;
wire net773;
wire net774_c1;
wire net774;
wire net775_c1;
wire net775;
wire net776_c1;
wire net776;
wire net777_c1;
wire net777;
wire net778_c1;
wire net778;
wire net779_c1;
wire net779;
wire net780_c1;
wire net780;
wire net781_c1;
wire net781;
wire net782_c1;
wire net782;
wire net783_c1;
wire net783;
wire net784_c1;
wire net784;
wire net785_c1;
wire net785;
wire net786_c1;
wire net786;
wire net787_c1;
wire net787;
wire net788_c1;
wire net788;
wire net789_c1;
wire net789;
wire net790_c1;
wire net790;
wire net791_c1;
wire net791;
wire net792_c1;
wire net792;
wire net793_c1;
wire net793;
wire net794_c1;
wire net794;
wire net795_c1;
wire net795;
wire net796_c1;
wire net796;
wire net797_c1;
wire net797;
wire net798_c1;
wire net798;
wire net799_c1;
wire net799;
wire net800_c1;
wire net800;
wire net801_c1;
wire net801;
wire net802_c1;
wire net802;
wire net803_c1;
wire net803;
wire net804_c1;
wire net804;
wire net805_c1;
wire net805;
wire net806_c1;
wire net806;
wire net807_c1;
wire net807;
wire net808_c1;
wire net808;
wire net809_c1;
wire net809;
wire net810_c1;
wire net810;
wire net811_c1;
wire net811;
wire net812_c1;
wire net812;
wire net813_c1;
wire net813;
wire net814_c1;
wire net814;
wire net815_c1;
wire net815;
wire net816_c1;
wire net816;
wire net817_c1;
wire net817;
wire net818_c1;
wire net818;
wire net819_c1;
wire net819;
wire net820_c1;
wire net820;
wire net821_c1;
wire net821;
wire net822_c1;
wire net822;
wire net823_c1;
wire net823;
wire net824_c1;
wire net824;
wire net825_c1;
wire net825;
wire net826_c1;
wire net826;
wire net827_c1;
wire net827;
wire net828_c1;
wire net828;
wire net829_c1;
wire net829;
wire net830_c1;
wire net830;
wire net831_c1;
wire net831;
wire net832_c1;
wire net832;
wire net833_c1;
wire net833;
wire net834_c1;
wire net834;
wire net835_c1;
wire net835;
wire net836_c1;
wire net836;
wire net837_c1;
wire net837;
wire net838_c1;
wire net838;
wire net839_c1;
wire net839;
wire net840_c1;
wire net840;
wire net841_c1;
wire net841;
wire net842_c1;
wire net842;
wire net843_c1;
wire net843;
wire net844_c1;
wire net844;
wire net845_c1;
wire net845;
wire net846_c1;
wire net846;
wire net847_c1;
wire net847;
wire net848_c1;
wire net848;
wire net849_c1;
wire net849;
wire net850_c1;
wire net850;
wire net851_c1;
wire net851;
wire net852_c1;
wire net852;
wire net853_c1;
wire net853;
wire net854_c1;
wire net854;
wire net855_c1;
wire net855;
wire net856_c1;
wire net856;
wire net857_c1;
wire net857;
wire net858_c1;
wire net858;
wire net859_c1;
wire net859;
wire net860_c1;
wire net860;
wire net861_c1;
wire net861;
wire net862_c1;
wire net862;
wire net863_c1;
wire net863;
wire net864_c1;
wire net864;
wire net865_c1;
wire net865;
wire net866_c1;
wire net866;
wire net867_c1;
wire net867;
wire net868_c1;
wire net868;
wire net869_c1;
wire net869;
wire net870_c1;
wire net870;
wire net871_c1;
wire net871;
wire net872_c1;
wire net872;
wire net873_c1;
wire net873;
wire net874_c1;
wire net874;
wire net875_c1;
wire net875;
wire net876_c1;
wire net876;
wire net877_c1;
wire net877;
wire net878_c1;
wire net878;
wire net879_c1;
wire net879;
wire net880_c1;
wire net880;
wire net881_c1;
wire net881;
wire net882_c1;
wire net882;
wire net883_c1;
wire net883;
wire net884_c1;
wire net884;
wire net885_c1;
wire net885;
wire net886_c1;
wire net886;
wire net887_c1;
wire net887;
wire net888_c1;
wire net888;
wire net889_c1;
wire net889;
wire net890_c1;
wire net890;
wire net891_c1;
wire net891;
wire net892_c1;
wire net892;
wire net893_c1;
wire net893;
wire net894_c1;
wire net894;
wire net895_c1;
wire net895;
wire net896_c1;
wire net896;
wire net897_c1;
wire net897;
wire net898_c1;
wire net898;
wire net899_c1;
wire net899;
wire net900_c1;
wire net900;
wire net901_c1;
wire net901;
wire net902_c1;
wire net902;
wire net903_c1;
wire net903;
wire net904_c1;
wire net904;
wire net905_c1;
wire net905;
wire net906_c1;
wire net906;
wire net907_c1;
wire net907;
wire net908_c1;
wire net908;
wire net909_c1;
wire net909;
wire net910_c1;
wire net910;
wire net911_c1;
wire net911;
wire net912_c1;
wire net912;
wire net913_c1;
wire net913;
wire net914_c1;
wire net914;
wire net915_c1;
wire net915;
wire net916_c1;
wire net916;
wire net917_c1;
wire net917;
wire net918_c1;
wire net918;
wire net919_c1;
wire net919;
wire net920_c1;
wire net920;
wire net921_c1;
wire net921;
wire net922_c1;
wire net922;
wire net923_c1;
wire net923;
wire net924_c1;
wire net924;
wire net925_c1;
wire net925;
wire net926_c1;
wire net926;
wire net927_c1;
wire net927;
wire net928_c1;
wire net928;
wire net929_c1;
wire net929;
wire net930_c1;
wire net930;
wire net931_c1;
wire net931;
wire net932_c1;
wire net932;
wire net933_c1;
wire net933;
wire net934_c1;
wire net934;
wire net935_c1;
wire net935;
wire net936_c1;
wire net936;
wire net937_c1;
wire net937;
wire net938_c1;
wire net938;
wire net939_c1;
wire net939;
wire net940_c1;
wire net940;
wire net941_c1;
wire net941;
wire net942_c1;
wire net942;
wire net943_c1;
wire net943;
wire net944_c1;
wire net944;
wire net945_c1;
wire net945;
wire net946_c1;
wire net946;
wire net947_c1;
wire net947;
wire net948_c1;
wire net948;
wire net949_c1;
wire net949;
wire net950_c1;
wire net950;
wire net951_c1;
wire net951;
wire net952_c1;
wire net952;
wire net953_c1;
wire net953;
wire net954_c1;
wire net954;
wire net955_c1;
wire net955;
wire net956_c1;
wire net956;
wire net957_c1;
wire net957;
wire net958_c1;
wire net958;
wire net959_c1;
wire net959;
wire net960_c1;
wire net960;
wire net961_c1;
wire net961;
wire net962_c1;
wire net962;
wire net963_c1;
wire net963;
wire net964_c1;
wire net964;
wire net965_c1;
wire net965;
wire net966_c1;
wire net966;
wire net967_c1;
wire net967;
wire net968_c1;
wire net968;
wire net969_c1;
wire net969;
wire net970_c1;
wire net970;
wire net971_c1;
wire net971;
wire net972_c1;
wire net972;
wire net973_c1;
wire net973;
wire net974_c1;
wire net974;
wire net975_c1;
wire net975;
wire net976_c1;
wire net976;
wire net977_c1;
wire net977;
wire net978_c1;
wire net978;
wire net979_c1;
wire net979;
wire net980_c1;
wire net980;
wire net981_c1;
wire net981;
wire net982_c1;
wire net982;
wire net983_c1;
wire net983;
wire net984_c1;
wire net984;
wire net985_c1;
wire net985;
wire net986_c1;
wire net986;
wire net987_c1;
wire net987;
wire net988_c1;
wire net988;
wire net989_c1;
wire net989;
wire net990_c1;
wire net990;
wire net991_c1;
wire net991;
wire net992_c1;
wire net992;
wire net993_c1;
wire net993;
wire net994_c1;
wire net994;
wire net995_c1;
wire net995;
wire net996_c1;
wire net996;
wire net997_c1;
wire net997;
wire net998_c1;
wire net998;
wire net999_c1;
wire net999;
wire net1000_c1;
wire net1000;
wire net1001_c1;
wire net1001;
wire net1002_c1;
wire net1002;
wire net1003_c1;
wire net1003;
wire net1004_c1;
wire net1004;
wire net1005_c1;
wire net1005;
wire net1006_c1;
wire net1006;
wire net1007_c1;
wire net1007;
wire net1008_c1;
wire net1008;
wire net1009_c1;
wire net1009;
wire net1010_c1;
wire net1010;
wire net1011_c1;
wire net1011;
wire net1012_c1;
wire net1012;
wire net1013_c1;
wire net1013;
wire net1014_c1;
wire net1014;
wire net1015_c1;
wire net1015;
wire net1016_c1;
wire net1016;
wire net1017_c1;
wire net1017;
wire net1018_c1;
wire net1018;
wire net1019_c1;
wire net1019;
wire net1020_c1;
wire net1020;
wire net1021_c1;
wire net1021;
wire net1022_c1;
wire net1022;
wire net1023_c1;
wire net1023;
wire net1024_c1;
wire net1024;
wire net1025_c1;
wire net1025;
wire net1026_c1;
wire net1026;
wire net1027_c1;
wire net1027;
wire net1028_c1;
wire net1028;
wire net1029_c1;
wire net1029;
wire net1030_c1;
wire net1030;
wire net1031_c1;
wire net1031;
wire net1032_c1;
wire net1032;
wire net1033_c1;
wire net1033;
wire net1034_c1;
wire net1034;
wire net1035_c1;
wire net1035;
wire net1036_c1;
wire net1036;
wire net1037_c1;
wire net1037;
wire net1038_c1;
wire net1038;
wire net1039_c1;
wire net1039;
wire net1040_c1;
wire net1040;
wire net1041_c1;
wire net1041;
wire net1042_c1;
wire net1042;
wire net1043_c1;
wire net1043;
wire net1044_c1;
wire net1044;
wire net1045_c1;
wire net1045;
wire net1046_c1;
wire net1046;
wire net1047_c1;
wire net1047;
wire net1048_c1;
wire net1048;
wire net1049_c1;
wire net1049;
wire net1050_c1;
wire net1050;
wire net1051_c1;
wire net1051;
wire net1052_c1;
wire net1052;
wire net1053_c1;
wire net1053;
wire net1054_c1;
wire net1054;
wire net1055_c1;
wire net1055;
wire net1056_c1;
wire net1056;
wire net1057_c1;
wire net1057;
wire net1058_c1;
wire net1058;
wire net1059_c1;
wire net1059;
wire net1060_c1;
wire net1060;
wire net1061_c1;
wire net1061;
wire net1062_c1;
wire net1062;
wire net1063_c1;
wire net1063;
wire net1064_c1;
wire net1064;
wire net1065_c1;
wire net1065;
wire net1066_c1;
wire net1066;
wire net1067_c1;
wire net1067;
wire net1068_c1;
wire net1068;
wire net1069_c1;
wire net1069;
wire net1070_c1;
wire net1070;
wire net1071_c1;
wire net1071;
wire net1072_c1;
wire net1072;
wire net1073_c1;
wire net1073;
wire net1074_c1;
wire net1074;
wire net1075_c1;
wire net1075;
wire net1076_c1;
wire net1076;
wire net1077_c1;
wire net1077;
wire net1078_c1;
wire net1078;
wire net1079_c1;
wire net1079;
wire net1080_c1;
wire net1080;
wire net1081_c1;
wire net1081;
wire net1082_c1;
wire net1082;
wire net1083_c1;
wire net1083;
wire net1084_c1;
wire net1084;
wire net1085_c1;
wire net1085;
wire net1086_c1;
wire net1086;
wire net1087_c1;
wire net1087;
wire net1088_c1;
wire net1088;
wire net1089_c1;
wire net1089;
wire net1090_c1;
wire net1090;
wire net1091_c1;
wire net1091;
wire net1092_c1;
wire net1092;
wire net1093_c1;
wire net1093;
wire net1094_c1;
wire net1094;
wire net1095_c1;
wire net1095;
wire net1096_c1;
wire net1096;
wire net1097_c1;
wire net1097;
wire net1098_c1;
wire net1098;
wire net1099_c1;
wire net1099;
wire net1100_c1;
wire net1100;
wire net1101_c1;
wire net1101;
wire net1102_c1;
wire net1102;
wire net1103_c1;
wire net1103;
wire net1104_c1;
wire net1104;
wire net1105_c1;
wire net1105;
wire net1106_c1;
wire net1106;
wire net1107_c1;
wire net1107;
wire net1108_c1;
wire net1108;
wire net1109_c1;
wire net1109;
wire net1110_c1;
wire net1110;
wire net1111_c1;
wire net1111;
wire net1112_c1;
wire net1112;
wire net1113_c1;
wire net1113;
wire net1114_c1;
wire net1114;
wire net1115_c1;
wire net1115;
wire net1116_c1;
wire net1116;
wire net1117_c1;
wire net1117;
wire net1118_c1;
wire net1118;
wire net1119_c1;
wire net1119;
wire net1120_c1;
wire net1120;
wire net1121_c1;
wire net1121;
wire net1122_c1;
wire net1122;
wire net1123_c1;
wire net1123;
wire net1124_c1;
wire net1124;
wire net1125_c1;
wire net1125;
wire net1126_c1;
wire net1126;
wire net1127_c1;
wire net1127;
wire net1128_c1;
wire net1128;
wire net1129_c1;
wire net1129;
wire net1130_c1;
wire net1130;
wire net1131_c1;
wire net1131;
wire net1132_c1;
wire net1132;
wire net1133_c1;
wire net1133;
wire net1134_c1;
wire net1134;
wire net1135_c1;
wire net1135;
wire net1136_c1;
wire net1136;
wire net1137_c1;
wire net1137;
wire net1138_c1;
wire net1138;
wire net1139_c1;
wire net1139;
wire net1140_c1;
wire net1140;
wire net1141_c1;
wire net1141;
wire net1142_c1;
wire net1142;
wire net1143_c1;
wire net1143;
wire net1144_c1;
wire net1144;
wire net1145_c1;
wire net1145;
wire net1146_c1;
wire net1146;
wire net1147_c1;
wire net1147;
wire net1148_c1;
wire net1148;
wire net1149_c1;
wire net1149;
wire net1150_c1;
wire net1150;
wire net1151_c1;
wire net1151;
wire net1152_c1;
wire net1152;
wire net1153_c1;
wire net1153;
wire net1154_c1;
wire net1154;
wire net1155_c1;
wire net1155;
wire net1156_c1;
wire net1156;
wire net1157_c1;
wire net1157;
wire net1158_c1;
wire net1158;
wire net1159_c1;
wire net1159;
wire net1160_c1;
wire net1160;
wire net1161_c1;
wire net1161;
wire net1162_c1;
wire net1162;
wire net1163_c1;
wire net1163;
wire net1164_c1;
wire net1164;
wire net1165_c1;
wire net1165;
wire net1166_c1;
wire net1166;
wire net1167_c1;
wire net1167;
wire net1168_c1;
wire net1168;
wire net1169_c1;
wire net1169;
wire net1170_c1;
wire net1170;
wire net1171_c1;
wire net1171;
wire net1172_c1;
wire net1172;
wire net1173_c1;
wire net1173;
wire net1174_c1;
wire net1174;
wire net1175_c1;
wire net1175;
wire net1176_c1;
wire net1176;
wire net1177_c1;
wire net1177;
wire net1178_c1;
wire net1178;
wire net1179_c1;
wire net1179;
wire net1180_c1;
wire net1180;
wire net1181_c1;
wire net1181;
wire net1182_c1;
wire net1182;
wire net1183_c1;
wire net1183;
wire net1184_c1;
wire net1184;
wire net1185_c1;
wire net1185;
wire net1186_c1;
wire net1186;
wire net1187_c1;
wire net1187;
wire net1188_c1;
wire net1188;
wire net1189_c1;
wire net1189;
wire net1190_c1;
wire net1190;
wire net1191_c1;
wire net1191;
wire net1192_c1;
wire net1192;
wire net1193_c1;
wire net1193;
wire net1194_c1;
wire net1194;
wire net1195_c1;
wire net1195;
wire net1196_c1;
wire net1196;
wire net1197_c1;
wire net1197;
wire net1198_c1;
wire net1198;
wire net1199_c1;
wire net1199;
wire net1200_c1;
wire net1200;
wire net1201_c1;
wire net1201;
wire net1202_c1;
wire net1202;
wire net1203_c1;
wire net1203;
wire net1204_c1;
wire net1204;
wire net1205_c1;
wire net1205;
wire net1206_c1;
wire net1206;
wire net1207_c1;
wire net1207;
wire net1208_c1;
wire net1208;
wire net1209_c1;
wire net1209;
wire net1210_c1;
wire net1210;
wire net1211_c1;
wire net1211;
wire net1212_c1;
wire net1212;
wire net1213_c1;
wire net1213;
wire net1214_c1;
wire net1214;
wire net1215_c1;
wire net1215;
wire net1216_c1;
wire net1216;
wire net1217_c1;
wire net1217;
wire net1218_c1;
wire net1218;
wire net1219_c1;
wire net1219;
wire net1220_c1;
wire net1220;
wire net1221_c1;
wire net1221;
wire net1222_c1;
wire net1222;
wire net1223_c1;
wire net1223;
wire net1224_c1;
wire net1224;
wire net1225_c1;
wire net1225;
wire net1226_c1;
wire net1226;
wire net1227_c1;
wire net1227;
wire net1228_c1;
wire net1228;
wire net1229_c1;
wire net1229;
wire net1230_c1;
wire net1230;
wire net1231_c1;
wire net1231;
wire net1232_c1;
wire net1232;
wire net1233_c1;
wire net1233;
wire net1234_c1;
wire net1234;
wire net1235_c1;
wire net1235;
wire net1236_c1;
wire net1236;
wire net1237_c1;
wire net1237;
wire net1238_c1;
wire net1238;
wire net1239_c1;
wire net1239;
wire net1240_c1;
wire net1240;
wire net1241_c1;
wire net1241;
wire net1242_c1;
wire net1242;
wire net1243_c1;
wire net1243;
wire net1244_c1;
wire net1244;
wire net1245_c1;
wire net1245;
wire net1246_c1;
wire net1246;
wire net1247_c1;
wire net1247;
wire net1248_c1;
wire net1248;
wire net1249_c1;
wire net1249;
wire net1250_c1;
wire net1250;
wire net1251_c1;
wire net1251;
wire net1252_c1;
wire net1252;
wire net1253_c1;
wire net1253;
wire net1254_c1;
wire net1254;
wire net1255_c1;
wire net1255;
wire net1256_c1;
wire net1256;
wire net1257_c1;
wire net1257;
wire net1258_c1;
wire net1258;
wire net1259_c1;
wire net1259;
wire net1260_c1;
wire net1260;
wire net1261_c1;
wire net1261;
wire net1262_c1;
wire net1262;
wire net1263_c1;
wire net1263;
wire net1264_c1;
wire net1264;
wire net1265_c1;
wire net1265;
wire net1266_c1;
wire net1266;
wire net1267_c1;
wire net1267;
wire net1268_c1;
wire net1268;
wire net1269_c1;
wire net1269;
wire net1270_c1;
wire net1270;
wire net1271_c1;
wire net1271;
wire net1272_c1;
wire net1272;
wire net1273_c1;
wire net1273;
wire net1274_c1;
wire net1274;
wire net1275_c1;
wire net1275;
wire net1276_c1;
wire net1276;
wire net1277_c1;
wire net1277;
wire net1278_c1;
wire net1278;
wire net1279_c1;
wire net1279;
wire net1280_c1;
wire net1280;
wire net1281_c1;
wire net1281;
wire net1282_c1;
wire net1282;
wire net1283_c1;
wire net1283;
wire net1284_c1;
wire net1284;
wire net1285_c1;
wire net1285;
wire net1286_c1;
wire net1286;
wire net1287_c1;
wire net1287;
wire net1288_c1;
wire net1288;
wire net1289_c1;
wire net1289;
wire net1290_c1;
wire net1290;
wire net1291_c1;
wire net1291;
wire net1292_c1;
wire net1292;
wire net1293_c1;
wire net1293;
wire net1294_c1;
wire net1294;
wire net1295_c1;
wire net1295;
wire net1296_c1;
wire net1296;
wire net1297_c1;
wire net1297;
wire net1298_c1;
wire net1298;
wire net1299_c1;
wire net1299;
wire net1300_c1;
wire net1300;
wire net1301_c1;
wire net1301;
wire net1302_c1;
wire net1302;
wire net1303_c1;
wire net1303;
wire net1304_c1;
wire net1304;
wire net1305_c1;
wire net1305;
wire net1306_c1;
wire net1306;
wire net1307_c1;
wire net1307;
wire net1308_c1;
wire net1308;
wire net1309_c1;
wire net1309;
wire net1310_c1;
wire net1310;
wire net1311_c1;
wire net1311;
wire net1312_c1;
wire net1312;
wire net1313_c1;
wire net1313;
wire net1314_c1;
wire net1314;
wire net1315_c1;
wire net1315;
wire net1316_c1;
wire net1316;
wire net1317_c1;
wire net1317;
wire net1318_c1;
wire net1318;
wire net1319_c1;
wire net1319;
wire net1320_c1;
wire net1320;
wire net1321_c1;
wire net1321;
wire net1322_c1;
wire net1322;
wire net1323_c1;
wire net1323;
wire net1324_c1;
wire net1324;
wire net1325_c1;
wire net1325;
wire net1326_c1;
wire net1326;
wire net1327_c1;
wire net1327;
wire net1328_c1;
wire net1328;
wire net1329_c1;
wire net1329;
wire net1330_c1;
wire net1330;
wire net1331_c1;
wire net1331;
wire net1332_c1;
wire net1332;
wire net1333_c1;
wire net1333;
wire net1334_c1;
wire net1334;
wire net1335_c1;
wire net1335;
wire net1336_c1;
wire net1336;
wire net1337_c1;
wire net1337;
wire net1338_c1;
wire net1338;
wire net1339_c1;
wire net1339;
wire net1340_c1;
wire net1340;
wire net1341_c1;
wire net1341;
wire net1342_c1;
wire net1342;
wire net1343_c1;
wire net1343;
wire net1344_c1;
wire net1344;
wire net1345_c1;
wire net1345;
wire net1346_c1;
wire net1346;
wire net1347_c1;
wire net1347;
wire net1348_c1;
wire net1348;
wire net1349_c1;
wire net1349;
wire net1350_c1;
wire net1350;
wire net1351_c1;
wire net1351;
wire net1352_c1;
wire net1352;
wire net1353_c1;
wire net1353;
wire net1354_c1;
wire net1354;
wire net1355_c1;
wire net1355;
wire net1356_c1;
wire net1356;
wire net1357_c1;
wire net1357;
wire net1358_c1;
wire net1358;
wire net1359_c1;
wire net1359;
wire net1360_c1;
wire net1360;
wire net1361_c1;
wire net1361;
wire net1362_c1;
wire net1362;
wire net1363_c1;
wire net1363;
wire net1364_c1;
wire net1364;
wire net1365_c1;
wire net1365;
wire net1366_c1;
wire net1366;
wire net1367_c1;
wire net1367;
wire net1368_c1;
wire net1368;
wire net1369_c1;
wire net1369;
wire net1370_c1;
wire net1370;
wire net1371_c1;
wire net1371;
wire net1372_c1;
wire net1372;
wire net1373_c1;
wire net1373;
wire net1374_c1;
wire net1374;
wire net1375_c1;
wire net1375;
wire net1376_c1;
wire net1376;
wire net1377_c1;
wire net1377;
wire net1378_c1;
wire net1378;
wire net1379_c1;
wire net1379;
wire net1380_c1;
wire net1380;
wire net1381_c1;
wire net1381;
wire net1382_c1;
wire net1382;
wire net1383_c1;
wire net1383;
wire net1384_c1;
wire net1384;
wire net1385_c1;
wire net1385;
wire net1386_c1;
wire net1386;
wire net1387_c1;
wire net1387;
wire net1388_c1;
wire net1388;
wire net1389_c1;
wire net1389;
wire net1390_c1;
wire net1390;
wire net1391_c1;
wire net1391;
wire net1392_c1;
wire net1392;
wire net1393_c1;
wire net1393;
wire net1394_c1;
wire net1394;
wire net1395_c1;
wire net1395;
wire net1396_c1;
wire net1396;
wire net1397_c1;
wire net1397;
wire net1398_c1;
wire net1398;
wire net1399_c1;
wire net1399;
wire net1400_c1;
wire net1400;
wire net1401_c1;
wire net1401;
wire net1402_c1;
wire net1402;
wire net1403_c1;
wire net1403;
wire net1404_c1;
wire net1404;
wire net1405_c1;
wire net1405;
wire net1406_c1;
wire net1406;
wire net1407_c1;
wire net1407;
wire net1408_c1;
wire net1408;
wire net1409_c1;
wire net1409;
wire net1410_c1;
wire net1410;
wire net1411_c1;
wire net1411;
wire net1412_c1;
wire net1412;
wire net1413_c1;
wire net1413;
wire net1414_c1;
wire net1414;
wire net1415_c1;
wire net1415;
wire net1416_c1;
wire net1416;
wire net1417_c1;
wire net1417;
wire net1418_c1;
wire net1418;
wire net1419_c1;
wire net1419;
wire net1420_c1;
wire net1420;
wire net1421_c1;
wire net1421;
wire net1422_c1;
wire net1422;
wire net1423_c1;
wire net1423;
wire net1424_c1;
wire net1424;
wire net1425_c1;
wire net1425;
wire net1426_c1;
wire net1426;
wire net1427_c1;
wire net1427;
wire net1428_c1;
wire net1428;
wire net1429_c1;
wire net1429;
wire net1430_c1;
wire net1430;
wire net1431_c1;
wire net1431;
wire net1432_c1;
wire net1432;
wire net1433_c1;
wire net1433;
wire net1434_c1;
wire net1434;
wire net1435_c1;
wire net1435;
wire net1436_c1;
wire net1436;
wire net1437_c1;
wire net1437;
wire net1438_c1;
wire net1438;
wire net1439_c1;
wire net1439;
wire net1440_c1;
wire net1440;
wire net1441_c1;
wire net1441;
wire net1442_c1;
wire net1442;
wire net1443_c1;
wire net1443;
wire net1444_c1;
wire net1444;
wire net1445_c1;
wire net1445;
wire net1446_c1;
wire net1446;
wire net1447_c1;
wire net1447;
wire net1448_c1;
wire net1448;
wire net1449_c1;
wire net1449;
wire net1450_c1;
wire net1450;
wire net1451_c1;
wire net1451;
wire net1452_c1;
wire net1452;
wire net1453_c1;
wire net1453;
wire net1454_c1;
wire net1454;
wire net1455_c1;
wire net1455;
wire net1456_c1;
wire net1456;
wire net1457_c1;
wire net1457;
wire net1458_c1;
wire net1458;
wire net1459_c1;
wire net1459;
wire net1460_c1;
wire net1460;
wire net1461_c1;
wire net1461;
wire net1462_c1;
wire net1462;
wire net1463_c1;
wire net1463;
wire net1464_c1;
wire net1464;
wire net1465_c1;
wire net1465;
wire net1466_c1;
wire net1466;
wire net1467_c1;
wire net1467;
wire net1468_c1;
wire net1468;
wire net1469_c1;
wire net1469;
wire net1470_c1;
wire net1470;
wire net1471_c1;
wire net1471;
wire net1472_c1;
wire net1472;
wire net1473_c1;
wire net1473;
wire net1474_c1;
wire net1474;
wire net1475_c1;
wire net1475;
wire net1476_c1;
wire net1476;
wire net1477_c1;
wire net1477;
wire net1478_c1;
wire net1478;
wire net1479_c1;
wire net1479;
wire net1480_c1;
wire net1480;
wire net1481_c1;
wire net1481;
wire net1482_c1;
wire net1482;
wire net1483_c1;
wire net1483;
wire net1484_c1;
wire net1484;
wire net1485_c1;
wire net1485;
wire net1486_c1;
wire net1486;
wire net1487_c1;
wire net1487;
wire net1488_c1;
wire net1488;
wire net1489_c1;
wire net1489;
wire net1490_c1;
wire net1490;
wire net1491_c1;
wire net1491;
wire net1492_c1;
wire net1492;
wire net1493_c1;
wire net1493;
wire net1494_c1;
wire net1494;
wire net1495_c1;
wire net1495;
wire net1496_c1;
wire net1496;
wire net1497_c1;
wire net1497;
wire net1498_c1;
wire net1498;
wire net1499_c1;
wire net1499;
wire net1500_c1;
wire net1500;
wire net1501_c1;
wire net1501;
wire net1502_c1;
wire net1502;
wire net1503_c1;
wire net1503;
wire net1504_c1;
wire net1504;
wire net1505_c1;
wire net1505;
wire net1506_c1;
wire net1506;
wire net1507_c1;
wire net1507;
wire net1508_c1;
wire net1508;
wire net1509_c1;
wire net1509;
wire net1510_c1;
wire net1510;
wire net1511_c1;
wire net1511;
wire net1512_c1;
wire net1512;
wire net1513_c1;
wire net1513;
wire net1514_c1;
wire net1514;
wire net1515_c1;
wire net1515;
wire net1516_c1;
wire net1516;
wire net1517_c1;
wire net1517;
wire net1518_c1;
wire net1518;
wire net1519_c1;
wire net1519;
wire net1520_c1;
wire net1520;
wire net1521_c1;
wire net1521;
wire net1522_c1;
wire net1522;
wire net1523_c1;
wire net1523;
wire net1524_c1;
wire net1524;
wire net1525_c1;
wire net1525;
wire net1526_c1;
wire net1526;
wire net1527_c1;
wire net1527;
wire net1528_c1;
wire net1528;
wire net1529_c1;
wire net1529;
wire net1530_c1;
wire net1530;
wire net1531_c1;
wire net1531;
wire net1532_c1;
wire net1532;
wire net1533_c1;
wire net1533;
wire net1534_c1;
wire net1534;
wire net1535_c1;
wire net1535;
wire net1536_c1;
wire net1536;
wire net1537_c1;
wire net1537;
wire net1538_c1;
wire net1538;
wire net1539_c1;
wire net1539;
wire net1540_c1;
wire net1540;
wire net1541_c1;
wire net1541;
wire net1542_c1;
wire net1542;
wire net1543_c1;
wire net1543;
wire net1544_c1;
wire net1544;
wire net1545_c1;
wire net1545;
wire net1546_c1;
wire net1546;
wire net1547_c1;
wire net1547;
wire net1548_c1;
wire net1548;
wire net1549_c1;
wire net1549;
wire net1550_c1;
wire net1550;
wire net1551_c1;
wire net1551;
wire net1552_c1;
wire net1552;
wire net1553_c1;
wire net1553;
wire net1554_c1;
wire net1554;
wire net1555_c1;
wire net1555;
wire net1556_c1;
wire net1556;
wire net1557_c1;
wire net1557;
wire net1558_c1;
wire net1558;
wire net1559_c1;
wire net1559;
wire net1560_c1;
wire net1560;
wire net1561_c1;
wire net1561;
wire net1562_c1;
wire net1562;
wire net1563_c1;
wire net1563;
wire net1564_c1;
wire net1564;
wire net1565_c1;
wire net1565;
wire net1566_c1;
wire net1566;
wire net1567_c1;
wire net1567;
wire net1568_c1;
wire net1568;
wire net1569_c1;
wire net1569;
wire net1570_c1;
wire net1570;
wire net1571_c1;
wire net1571;
wire net1572_c1;
wire net1572;
wire net1573_c1;
wire net1573;
wire net1574_c1;
wire net1574;
wire net1575_c1;
wire net1575;
wire net1576_c1;
wire net1576;
wire net1577_c1;
wire net1577;
wire net1578_c1;
wire net1578;
wire net1579_c1;
wire net1579;
wire net1580_c1;
wire net1580;
wire net1581_c1;
wire net1581;
wire net1582_c1;
wire net1582;
wire net1583_c1;
wire net1583;
wire net1584_c1;
wire net1584;
wire net1585_c1;
wire net1585;
wire net1586_c1;
wire net1586;
wire net1587_c1;
wire net1587;
wire net1588_c1;
wire net1588;
wire net1589_c1;
wire net1589;
wire net1590_c1;
wire net1590;
wire net1591_c1;
wire net1591;
wire net1592_c1;
wire net1592;
wire net1593_c1;
wire net1593;
wire net1594_c1;
wire net1594;
wire net1595_c1;
wire net1595;
wire net1596_c1;
wire net1596;
wire net1597_c1;
wire net1597;
wire net1598_c1;
wire net1598;
wire net1599_c1;
wire net1599;
wire net1600_c1;
wire net1600;
wire net1601_c1;
wire net1601;
wire net1602_c1;
wire net1602;
wire net1603_c1;
wire net1603;
wire net1604_c1;
wire net1604;
wire net1605_c1;
wire net1605;
wire net1606_c1;
wire net1606;
wire net1607_c1;
wire net1607;
wire net1608_c1;
wire net1608;
wire net1609_c1;
wire net1609;
wire net1610_c1;
wire net1610;
wire net1611_c1;
wire net1611;
wire net1612_c1;
wire net1612;
wire net1613_c1;
wire net1613;
wire net1614_c1;
wire net1614;
wire net1615_c1;
wire net1615;
wire net1616_c1;
wire net1616;
wire net1617_c1;
wire net1617;
wire net1618_c1;
wire net1618;
wire net1619_c1;
wire net1619;
wire net1620_c1;
wire net1620;
wire net1621_c1;
wire net1621;
wire net1622_c1;
wire net1622;
wire net1623_c1;
wire net1623;
wire net1624_c1;
wire net1624;
wire net1625_c1;
wire net1625;
wire net1626_c1;
wire net1626;
wire net1627_c1;
wire net1627;
wire net1628_c1;
wire net1628;
wire net1629_c1;
wire net1629;
wire net1630_c1;
wire net1630;
wire net1631_c1;
wire net1631;
wire net1632_c1;
wire net1632;
wire net1633_c1;
wire net1633;
wire net1634_c1;
wire net1634;
wire net1635_c1;
wire net1635;
wire net1636_c1;
wire net1636;
wire net1637_c1;
wire net1637;
wire net1638_c1;
wire net1638;
wire net1639_c1;
wire net1639;
wire net1640_c1;
wire net1640;
wire net1641_c1;
wire net1641;
wire net1642_c1;
wire net1642;
wire net1643_c1;
wire net1643;
wire net1644_c1;
wire net1644;
wire net1645_c1;
wire net1645;
wire net1646_c1;
wire net1646;
wire net1647_c1;
wire net1647;
wire net1648_c1;
wire net1648;
wire net1649_c1;
wire net1649;
wire net1650_c1;
wire net1650;
wire net1651_c1;
wire net1651;
wire net1652_c1;
wire net1652;
wire net1653_c1;
wire net1653;
wire net1654_c1;
wire net1654;
wire net1655_c1;
wire net1655;
wire net1656_c1;
wire net1656;
wire net1657_c1;
wire net1657;
wire net1658_c1;
wire net1658;
wire net1659_c1;
wire net1659;
wire net1660_c1;
wire net1660;
wire net1661_c1;
wire net1661;
wire net1662_c1;
wire net1662;
wire net1663_c1;
wire net1663;
wire net1664_c1;
wire net1664;
wire net1665_c1;
wire net1665;
wire net1666_c1;
wire net1666;
wire net1667_c1;
wire net1667;
wire net1668_c1;
wire net1668;
wire net1669_c1;
wire net1669;
wire net1670_c1;
wire net1670;
wire net1671_c1;
wire net1671;
wire net1672_c1;
wire net1672;
wire net1673_c1;
wire net1673;
wire net1674_c1;
wire net1674;
wire net1675_c1;
wire net1675;
wire net1676_c1;
wire net1676;
wire net1677_c1;
wire net1677;
wire net1678_c1;
wire net1678;
wire net1679_c1;
wire net1679;
wire net1680_c1;
wire net1680;
wire net1681_c1;
wire net1681;
wire net1682_c1;
wire net1682;
wire net1683_c1;
wire net1683;
wire net1684_c1;
wire net1684;
wire net1685_c1;
wire net1685;
wire net1686_c1;
wire net1686;
wire net1687_c1;
wire net1687;
wire net1688_c1;
wire net1688;
wire net1689_c1;
wire net1689;
wire net1690_c1;
wire net1690;
wire net1691_c1;
wire net1691;
wire net1692_c1;
wire net1692;
wire net1693_c1;
wire net1693;
wire net1694_c1;
wire net1694;
wire net1695_c1;
wire net1695;
wire net1696_c1;
wire net1696;
wire net1697_c1;
wire net1697;
wire net1698_c1;
wire net1698;
wire net1699_c1;
wire net1699;
wire net1700_c1;
wire net1700;
wire net1701_c1;
wire net1701;
wire net1702_c1;
wire net1702;
wire net1703_c1;
wire net1703;
wire net1704_c1;
wire net1704;
wire net1705_c1;
wire net1705;
wire net1706_c1;
wire net1706;
wire net1707_c1;
wire net1707;
wire net1708_c1;
wire net1708;
wire net1709_c1;
wire net1709;
wire net1710_c1;
wire net1710;
wire net1711_c1;
wire net1711;
wire net1712_c1;
wire net1712;
wire net1713_c1;
wire net1713;
wire net1714_c1;
wire net1714;
wire net1715_c1;
wire net1715;
wire net1716_c1;
wire net1716;
wire net1717_c1;
wire net1717;
wire net1718_c1;
wire net1718;
wire net1719_c1;
wire net1719;
wire net1720_c1;
wire net1720;
wire net1721_c1;
wire net1721;
wire net1722_c1;
wire net1722;
wire net1723_c1;
wire net1723;
wire net1724_c1;
wire net1724;
wire net1725_c1;
wire net1725;
wire net1726_c1;
wire net1726;
wire net1727_c1;
wire net1727;
wire net1728_c1;
wire net1728;
wire net1729_c1;
wire net1729;
wire net1730_c1;
wire net1730;
wire net1731_c1;
wire net1731;
wire net1732_c1;
wire net1732;
wire net1733_c1;
wire net1733;
wire net1734_c1;
wire net1734;
wire net1735_c1;
wire net1735;
wire net1736_c1;
wire net1736;
wire net1737_c1;
wire net1737;
wire net1738_c1;
wire net1738;
wire net1739_c1;
wire net1739;
wire net1740_c1;
wire net1740;
wire net1741_c1;
wire net1741;
wire net1742_c1;
wire net1742;
wire net1743_c1;
wire net1743;
wire net1744_c1;
wire net1744;
wire net1745_c1;
wire net1745;
wire net1746_c1;
wire net1746;
wire net1747_c1;
wire net1747;
wire net1748_c1;
wire net1748;
wire net1749_c1;
wire net1749;
wire net1750_c1;
wire net1750;
wire net1751_c1;
wire net1751;
wire net1752_c1;
wire net1752;
wire net1753_c1;
wire net1753;
wire net1754_c1;
wire net1754;
wire net1755_c1;
wire net1755;
wire net1756_c1;
wire net1756;
wire net1757_c1;
wire net1757;
wire net1758_c1;
wire net1758;
wire net1759_c1;
wire net1759;
wire net1760_c1;
wire net1760;
wire net1761_c1;
wire net1761;
wire net1762_c1;
wire net1762;
wire net1763_c1;
wire net1763;
wire net1764_c1;
wire net1764;
wire net1765_c1;
wire net1765;
wire net1766_c1;
wire net1766;
wire net1767_c1;
wire net1767;
wire net1768_c1;
wire net1768;
wire net1769_c1;
wire net1769;
wire net1770_c1;
wire net1770;
wire net1771_c1;
wire net1771;
wire net1772_c1;
wire net1772;
wire net1773_c1;
wire net1773;
wire net1774_c1;
wire net1774;
wire net1775_c1;
wire net1775;
wire net1776_c1;
wire net1776;
wire net1777_c1;
wire net1777;
wire net1778_c1;
wire net1778;
wire net1779_c1;
wire net1779;
wire net1780_c1;
wire net1780;
wire net1781_c1;
wire net1781;
wire net1782_c1;
wire net1782;
wire net1783_c1;
wire net1783;
wire net1784_c1;
wire net1784;
wire net1785_c1;
wire net1785;
wire net1786_c1;
wire net1786;
wire net1787_c1;
wire net1787;
wire net1788_c1;
wire net1788;
wire net1789_c1;
wire net1789;
wire net1790_c1;
wire net1790;
wire net1791_c1;
wire net1791;
wire net1792_c1;
wire net1792;
wire net1793_c1;
wire net1793;
wire net1794_c1;
wire net1794;
wire net1795_c1;
wire net1795;
wire net1796_c1;
wire net1796;
wire net1797_c1;
wire net1797;
wire net1798_c1;
wire net1798;
wire net1799_c1;
wire net1799;
wire net1800_c1;
wire net1800;
wire net1801_c1;
wire net1801;
wire net1802_c1;
wire net1802;
wire net1803_c1;
wire net1803;
wire net1804_c1;
wire net1804;
wire net1805_c1;
wire net1805;
wire net1806_c1;
wire net1806;
wire net1807_c1;
wire net1807;
wire net1808_c1;
wire net1808;
wire net1809_c1;
wire net1809;
wire net1810_c1;
wire net1810;
wire net1811_c1;
wire net1811;
wire net1812_c1;
wire net1812;
wire net1813_c1;
wire net1813;
wire net1814_c1;
wire net1814;
wire net1815_c1;
wire net1815;
wire net1816_c1;
wire net1816;
wire net1817_c1;
wire net1817;
wire net1818_c1;
wire net1818;
wire net1819_c1;
wire net1819;
wire net1820_c1;
wire net1820;
wire net1821_c1;
wire net1821;
wire net1822_c1;
wire net1822;
wire net1823_c1;
wire net1823;
wire net1824_c1;
wire net1824;
wire net1825_c1;
wire net1825;
wire net1826_c1;
wire net1826;
wire net1827_c1;
wire net1827;
wire net1828_c1;
wire net1828;
wire net1829_c1;
wire net1829;
wire net1830_c1;
wire net1830;
wire net1831_c1;
wire net1831;
wire net1832_c1;
wire net1832;
wire net1833_c1;
wire net1833;
wire net1834_c1;
wire net1834;
wire net1835_c1;
wire net1835;
wire net1836_c1;
wire net1836;
wire net1837_c1;
wire net1837;
wire net1838_c1;
wire net1838;
wire net1839_c1;
wire net1839;
wire net1840_c1;
wire net1840;
wire net1841_c1;
wire net1841;
wire net1842_c1;
wire net1842;
wire net1843_c1;
wire net1843;
wire net1844_c1;
wire net1844;
wire net1845_c1;
wire net1845;
wire net1846_c1;
wire net1846;
wire net1847_c1;
wire net1847;
wire net1848_c1;
wire net1848;
wire net1849_c1;
wire net1849;
wire net1850_c1;
wire net1850;
wire net1851_c1;
wire net1851;
wire net1852_c1;
wire net1852;
wire net1853_c1;
wire net1853;
wire net1854_c1;
wire net1854;
wire net1855_c1;
wire net1855;
wire net1856_c1;
wire net1856;
wire net1857_c1;
wire net1857;
wire net1858_c1;
wire net1858;
wire net1859_c1;
wire net1859;
wire net1860_c1;
wire net1860;
wire net1861_c1;
wire net1861;
wire net1862_c1;
wire net1862;
wire net1863_c1;
wire net1863;
wire net1864_c1;
wire net1864;
wire net1865_c1;
wire net1865;
wire net1866_c1;
wire net1866;
wire net1867_c1;
wire net1867;
wire net1868_c1;
wire net1868;
wire net1869_c1;
wire net1869;
wire net1870_c1;
wire net1870;
wire net1871_c1;
wire net1871;
wire net1872_c1;
wire net1872;
wire net1873_c1;
wire net1873;
wire net1874_c1;
wire net1874;
wire net1875_c1;
wire net1875;
wire net1876_c1;
wire net1876;
wire net1877_c1;
wire net1877;
wire net1878_c1;
wire net1878;
wire net1879_c1;
wire net1879;
wire net1880_c1;
wire net1880;
wire net1881_c1;
wire net1881;
wire net1882_c1;
wire net1882;
wire net1883_c1;
wire net1883;
wire net1884_c1;
wire net1884;
wire net1885_c1;
wire net1885;
wire net1886_c1;
wire net1886;
wire net1887_c1;
wire net1887;
wire net1888_c1;
wire net1888;
wire net1889_c1;
wire net1889;
wire net1890_c1;
wire net1890;
wire net1891_c1;
wire net1891;
wire net1892_c1;
wire net1892;
wire net1893_c1;
wire net1893;
wire net1894_c1;
wire net1894;
wire net1895_c1;
wire net1895;
wire net1896_c1;
wire net1896;
wire net1897_c1;
wire net1897;
wire net1898_c1;
wire net1898;
wire net1899_c1;
wire net1899;
wire net1900_c1;
wire net1900;
wire net1901_c1;
wire net1901;
wire net1902_c1;
wire net1902;
wire net1903_c1;
wire net1903;
wire net1904_c1;
wire net1904;
wire net1905_c1;
wire net1905;
wire net1906_c1;
wire net1906;
wire net1907_c1;
wire net1907;
wire net1908_c1;
wire net1908;
wire net1909_c1;
wire net1909;
wire net1910_c1;
wire net1910;
wire net1911_c1;
wire net1911;
wire net1912_c1;
wire net1912;
wire net1913_c1;
wire net1913;
wire net1914_c1;
wire net1914;
wire net1915_c1;
wire net1915;
wire net1916_c1;
wire net1916;
wire net1917_c1;
wire net1917;
wire net1918_c1;
wire net1918;
wire net1919_c1;
wire net1919;
wire net1920_c1;
wire net1920;
wire net1921_c1;
wire net1921;
wire net1922_c1;
wire net1922;
wire net1923_c1;
wire net1923;
wire net1924_c1;
wire net1924;
wire net1925_c1;
wire net1925;
wire net1926_c1;
wire net1926;
wire net1927_c1;
wire net1927;
wire net1928_c1;
wire net1928;
wire net1929_c1;
wire net1929;
wire net1930_c1;
wire net1930;
wire net1931_c1;
wire net1931;
wire net1932_c1;
wire net1932;
wire net1933_c1;
wire net1933;
wire net1934_c1;
wire net1934;
wire net1935_c1;
wire net1935;
wire net1936_c1;
wire net1936;
wire net1937_c1;
wire net1937;
wire net1938_c1;
wire net1938;
wire net1939_c1;
wire net1939;
wire net1940_c1;
wire net1940;
wire net1941_c1;
wire net1941;
wire net1942_c1;
wire net1942;
wire net1943_c1;
wire net1943;
wire net1944_c1;
wire net1944;
wire net1945_c1;
wire net1945;
wire net1946_c1;
wire net1946;
wire net1947_c1;
wire net1947;
wire net1948_c1;
wire net1948;
wire net1949_c1;
wire net1949;
wire net1950_c1;
wire net1950;
wire net1951_c1;
wire net1951;
wire net1952_c1;
wire net1952;
wire net1953_c1;
wire net1953;
wire net1954_c1;
wire net1954;
wire net1955_c1;
wire net1955;
wire net1956_c1;
wire net1956;
wire net1957_c1;
wire net1957;
wire net1958_c1;
wire net1958;
wire net1959_c1;
wire net1959;
wire net1960_c1;
wire net1960;
wire net1961_c1;
wire net1961;
wire net1962_c1;
wire net1962;
wire net1963_c1;
wire net1963;
wire net1964_c1;
wire net1964;
wire net1965_c1;
wire net1965;
wire net1966_c1;
wire net1966;
wire net1967_c1;
wire net1967;
wire net1968_c1;
wire net1968;
wire net1969_c1;
wire net1969;
wire net1970_c1;
wire net1970;
wire net1971_c1;
wire net1971;
wire net1972_c1;
wire net1972;
wire net1973_c1;
wire net1973;
wire net1974_c1;
wire net1974;
wire net1975_c1;
wire net1975;
wire net1976_c1;
wire net1976;
wire net1977_c1;
wire net1977;
wire net1978_c1;
wire net1978;
wire net1979_c1;
wire net1979;
wire net1980_c1;
wire net1980;
wire net1981_c1;
wire net1981;
wire net1982_c1;
wire net1982;
wire net1983_c1;
wire net1983;
wire net1984_c1;
wire net1984;
wire net1985_c1;
wire net1985;
wire net1986_c1;
wire net1986;
wire net1987_c1;
wire net1987;
wire net1988_c1;
wire net1988;
wire net1989_c1;
wire net1989;
wire net1990_c1;
wire net1990;
wire net1991_c1;
wire net1991;
wire net1992_c1;
wire net1992;
wire net1993_c1;
wire net1993;
wire net1994_c1;
wire net1994;
wire net1995_c1;
wire net1995;
wire net1996_c1;
wire net1996;
wire net1997_c1;
wire net1997;
wire net1998_c1;
wire net1998;
wire net1999_c1;
wire net1999;
wire net2000_c1;
wire net2000;
wire net2001_c1;
wire net2001;
wire net2002_c1;
wire net2002;
wire net2003_c1;
wire net2003;
wire net2004_c1;
wire net2004;
wire net2005_c1;
wire net2005;
wire net2006_c1;
wire net2006;
wire net2007_c1;
wire net2007;
wire net2008_c1;
wire net2008;
wire net2009_c1;
wire net2009;
wire net2010_c1;
wire net2010;
wire net2011_c1;
wire net2011;
wire net2012_c1;
wire net2012;
wire net2013_c1;
wire net2013;
wire net2014_c1;
wire net2014;
wire net2015_c1;
wire net2015;
wire net2016_c1;
wire net2016;
wire net2017_c1;
wire net2017;
wire net2018_c1;
wire net2018;
wire net2019_c1;
wire net2019;
wire net2020_c1;
wire net2020;
wire net2021_c1;
wire net2021;
wire net2022_c1;
wire net2022;
wire net2023_c1;
wire net2023;
wire net2024_c1;
wire net2024;
wire net2025_c1;
wire net2025;
wire net2026_c1;
wire net2026;
wire net2027_c1;
wire net2027;
wire net2028_c1;
wire net2028;
wire net2029_c1;
wire net2029;
wire net2030_c1;
wire net2030;
wire net2031_c1;
wire net2031;
wire net2032_c1;
wire net2032;
wire net2033_c1;
wire net2033;
wire net2034_c1;
wire net2034;
wire net2035_c1;
wire net2035;
wire net2036_c1;
wire net2036;
wire net2037_c1;
wire net2037;
wire net2038_c1;
wire net2038;
wire net2039_c1;
wire net2039;
wire net2040_c1;
wire net2040;
wire net2041_c1;
wire net2041;
wire net2042_c1;
wire net2042;
wire net2043_c1;
wire net2043;
wire net2044_c1;
wire net2044;
wire net2045_c1;
wire net2045;
wire net2046_c1;
wire net2046;
wire net2047_c1;
wire net2047;
wire net2048_c1;
wire net2048;
wire net2049_c1;
wire net2049;
wire net2050_c1;
wire net2050;
wire net2051_c1;
wire net2051;
wire net2052_c1;
wire net2052;
wire net2053_c1;
wire net2053;
wire net2054_c1;
wire net2054;
wire net2055_c1;
wire net2055;
wire net2056_c1;
wire net2056;
wire net2057_c1;
wire net2057;
wire net2058_c1;
wire net2058;
wire net2059_c1;
wire net2059;
wire net2060_c1;
wire net2060;
wire net2061_c1;
wire net2061;
wire net2062_c1;
wire net2062;
wire net2063_c1;
wire net2063;
wire net2064_c1;
wire net2064;
wire net2065_c1;
wire net2065;
wire net2066_c1;
wire net2066;
wire net2067_c1;
wire net2067;
wire net2068_c1;
wire net2068;
wire net2069_c1;
wire net2069;
wire net2070_c1;
wire net2070;
wire net2071_c1;
wire net2071;
wire net2072_c1;
wire net2072;
wire net2073_c1;
wire net2073;
wire net2074_c1;
wire net2074;
wire net2075_c1;
wire net2075;
wire net2076_c1;
wire net2076;
wire net2077_c1;
wire net2077;
wire net2078_c1;
wire net2078;
wire net2079_c1;
wire net2079;
wire net2080_c1;
wire net2080;
wire net2081_c1;
wire net2081;
wire net2082_c1;
wire net2082;
wire net2083_c1;
wire net2083;
wire net2084_c1;
wire net2084;
wire net2085_c1;
wire net2085;
wire net2086_c1;
wire net2086;
wire net2087_c1;
wire net2087;
wire net2088_c1;
wire net2088;
wire net2089_c1;
wire net2089;
wire net2090_c1;
wire net2090;
wire net2091_c1;
wire net2091;
wire net2092_c1;
wire net2092;
wire net2093_c1;
wire net2093;
wire net2094_c1;
wire net2094;
wire net2095_c1;
wire net2095;
wire net2096_c1;
wire net2096;
wire net2097_c1;
wire net2097;
wire net2098_c1;
wire net2098;
wire net2099_c1;
wire net2099;
wire net2100_c1;
wire net2100;
wire net2101_c1;
wire net2101;
wire net2102_c1;
wire net2102;
wire net2103_c1;
wire net2103;
wire net2104_c1;
wire net2104;
wire net2105_c1;
wire net2105;
wire net2106_c1;
wire net2106;
wire net2107_c1;
wire net2107;
wire net2108_c1;
wire net2108;
wire net2109_c1;
wire net2109;
wire net2110_c1;
wire net2110;
wire net2111_c1;
wire net2111;
wire net2112_c1;
wire net2112;
wire net2113_c1;
wire net2113;
wire net2114_c1;
wire net2114;
wire net2115_c1;
wire net2115;
wire net2116_c1;
wire net2116;
wire net2117_c1;
wire net2117;
wire net2118_c1;
wire net2118;
wire net2119_c1;
wire net2119;
wire net2120_c1;
wire net2120;
wire net2121_c1;
wire net2121;
wire net2122_c1;
wire net2122;
wire net2123_c1;
wire net2123;
wire net2124_c1;
wire net2124;
wire net2125_c1;
wire net2125;
wire net2126_c1;
wire net2126;
wire net2127_c1;
wire net2127;
wire net2128_c1;
wire net2128;
wire net2129_c1;
wire net2129;
wire net2130_c1;
wire net2130;
wire net2131_c1;
wire net2131;
wire net2132_c1;
wire net2132;
wire net2133_c1;
wire net2133;
wire net2134_c1;
wire net2134;
wire net2135_c1;
wire net2135;
wire net2136_c1;
wire net2136;
wire net2137_c1;
wire net2137;
wire net2138_c1;
wire net2138;
wire net2139_c1;
wire net2139;
wire net2140_c1;
wire net2140;
wire net2141_c1;
wire net2141;
wire net2142_c1;
wire net2142;
wire net2143_c1;
wire net2143;
wire net2144_c1;
wire net2144;
wire net2145_c1;
wire net2145;
wire net2146_c1;
wire net2146;
wire net2147_c1;
wire net2147;
wire net2148_c1;
wire net2148;
wire net2149_c1;
wire net2149;
wire net2150_c1;
wire net2150;
wire net2151_c1;
wire net2151;
wire net2152_c1;
wire net2152;
wire net2153_c1;
wire net2153;
wire net2154_c1;
wire net2154;
wire net2155_c1;
wire net2155;
wire net2156_c1;
wire net2156;
wire net2157_c1;
wire net2157;
wire net2158_c1;
wire net2158;
wire net2159_c1;
wire net2159;
wire net2160_c1;
wire net2160;
wire net2161_c1;
wire net2161;
wire net2162_c1;
wire net2162;
wire net2163_c1;
wire net2163;
wire net2164_c1;
wire net2164;
wire net2165_c1;
wire net2165;
wire net2166_c1;
wire net2166;
wire net2167_c1;
wire net2167;
wire net2168_c1;
wire net2168;
wire net2169_c1;
wire net2169;
wire net2170_c1;
wire net2170;
wire net2171_c1;
wire net2171;
wire net2172_c1;
wire net2172;
wire net2173_c1;
wire net2173;
wire net2174_c1;
wire net2174;
wire net2175_c1;
wire net2175;
wire net2176_c1;
wire net2176;
wire net2177_c1;
wire net2177;
wire net2178_c1;
wire net2178;
wire net2179_c1;
wire net2179;
wire net2180_c1;
wire net2180;
wire net2181_c1;
wire net2181;
wire net2182_c1;
wire net2182;
wire net2183_c1;
wire net2183;
wire net2184_c1;
wire net2184;
wire net2185_c1;
wire net2185;
wire net2186_c1;
wire net2186;
wire net2187_c1;
wire net2187;
wire net2188_c1;
wire net2188;
wire net2189_c1;
wire net2189;
wire net2190_c1;
wire net2190;
wire net2191_c1;
wire net2191;
wire net2192_c1;
wire net2192;
wire net2193_c1;
wire net2193;
wire net2194_c1;
wire net2194;
wire net2195_c1;
wire net2195;
wire net2196_c1;
wire net2196;
wire net2197_c1;
wire net2197;
wire net2198_c1;
wire net2198;
wire net2199_c1;
wire net2199;
wire net2200_c1;
wire net2200;
wire net2201_c1;
wire net2201;
wire net2202_c1;
wire net2202;
wire net2203_c1;
wire net2203;
wire net2204_c1;
wire net2204;
wire net2205_c1;
wire net2205;
wire net2206_c1;
wire net2206;
wire net2207_c1;
wire net2207;
wire net2208_c1;
wire net2208;
wire net2209_c1;
wire net2209;
wire net2210_c1;
wire net2210;
wire net2211_c1;
wire net2211;
wire net2212_c1;
wire net2212;
wire net2213_c1;
wire net2213;
wire net2214_c1;
wire net2214;
wire net2215_c1;
wire net2215;
wire net2216_c1;
wire net2216;
wire net2217_c1;
wire net2217;
wire net2218_c1;
wire net2218;
wire net2219_c1;
wire net2219;
wire net2220_c1;
wire net2220;
wire net2221_c1;
wire net2221;
wire net2222_c1;
wire net2222;
wire net2223_c1;
wire net2223;
wire net2224_c1;
wire net2224;
wire net2225_c1;
wire net2225;
wire net2226_c1;
wire net2226;
wire net2227_c1;
wire net2227;
wire net2228_c1;
wire net2228;
wire net2229_c1;
wire net2229;
wire net2230_c1;
wire net2230;
wire net2231_c1;
wire net2231;
wire net2232_c1;
wire net2232;
wire net2233_c1;
wire net2233;
wire net2234_c1;
wire net2234;
wire net2235_c1;
wire net2235;
wire net2236_c1;
wire net2236;
wire net2237_c1;
wire net2237;
wire net2238_c1;
wire net2238;
wire net2239_c1;
wire net2239;
wire net2240_c1;
wire net2240;
wire net2241_c1;
wire net2241;
wire net2242_c1;
wire net2242;
wire net2243_c1;
wire net2243;
wire net2244_c1;
wire net2244;
wire net2245_c1;
wire net2245;
wire net2246_c1;
wire net2246;
wire net2247_c1;
wire net2247;
wire net2248_c1;
wire net2248;
wire net2249_c1;
wire net2249;
wire net2250_c1;
wire net2250;
wire net2251_c1;
wire net2251;
wire net2252_c1;
wire net2252;
wire net2253_c1;
wire net2253;
wire net2254_c1;
wire net2254;
wire net2255_c1;
wire net2255;
wire net2256_c1;
wire net2256;
wire net2257_c1;
wire net2257;
wire net2258_c1;
wire net2258;
wire net2259_c1;
wire net2259;
wire net2260_c1;
wire net2260;
wire net2261_c1;
wire net2261;
wire net2262_c1;
wire net2262;
wire net2263_c1;
wire net2263;
wire net2264_c1;
wire net2264;
wire net2265_c1;
wire net2265;
wire net2266_c1;
wire net2266;
wire net2267_c1;
wire net2267;
wire net2268_c1;
wire net2268;
wire net2269_c1;
wire net2269;
wire net2270_c1;
wire net2270;
wire net2271_c1;
wire net2271;
wire net2272_c1;
wire net2272;
wire net2273_c1;
wire net2273;
wire net2274_c1;
wire net2274;
wire net2275_c1;
wire net2275;
wire net2276_c1;
wire net2276;
wire net2277_c1;
wire net2277;
wire net2278_c1;
wire net2278;
wire net2279_c1;
wire net2279;
wire net2280_c1;
wire net2280;
wire net2281_c1;
wire net2281;
wire net2282_c1;
wire net2282;
wire net2283_c1;
wire net2283;
wire GCLK_Pad;
wire net2284;
wire net2285_c1;
wire net2285;
wire net2286_c1;
wire net2286;
wire net2287_c1;
wire net2287;
wire net2288_c1;
wire net2288;
wire net2289_c1;
wire net2289;
wire net2290_c1;
wire net2290;
wire net2291_c1;
wire net2291;
wire net2292_c1;
wire net2292;
wire net2293_c1;
wire net2293;
wire net2294_c1;
wire net2294;
wire net2295_c1;
wire net2295;
wire net2296_c1;
wire net2296;
wire net2297_c1;
wire net2297;
wire net2298_c1;
wire net2298;
wire net2299_c1;
wire net2299;
wire net2300_c1;
wire net2300;
wire net2301_c1;
wire net2301;
wire net2302_c1;
wire net2302;
wire net2303_c1;
wire net2303;

DFFT DFFT_535__FPB_n1715(net1239,net563,net583_c1);
DFFT DFFT_471__FPB_n1651(net1238,net565,net584_c1);
DFFT DFFT_463__FPB_n1643(net2218,net566,net585_c1);
DFFT DFFT_455__FPB_n1635(net1237,net567,net586_c1);
DFFT DFFT_447__FPB_n1627(net1236,net568,net587_c1);
DFFT DFFT_439__FPB_n1619(net1235,net569,net588_c1);
DFFT DFFT_391__FPB_n1571(net1436,net570,net589_c1);
DFFT DFFT_383__FPB_n1563(net1234,net202,net590_c1);
DFFT DFFT_375__FPB_n1555(net1233,net571,net591_c1);
DFFT DFFT_367__FPB_n1547(net1232,net112,net600_c1);
DFFT DFFT_359__FPB_n1539(net1231,net102,net592_c1);
DFFT DFFT_295__FPB_n1475(net1230,net573,net601_c1);
DFFT DFFT_287__FPB_n1467(net1229,net574,net595_c1);
DFFT DFFT_279__FPB_n1459(net1228,net575,net596_c1);
DFFT DFFT_199__FPB_n1379(net1227,net577,net599_c1);
DFFT DFFT_519__FPB_n1699(net1226,net730,net731_c1);
DFFT DFFT_536__FPB_n1716(net1225,net583,net602_c1);
DFFT DFFT_528__FPB_n1708(net1224,net141,net603_c1);
DFFT DFFT_480__FPB_n1660(net1223,net700,net604_c1);
DFFT DFFT_472__FPB_n1652(net1222,net584,net605_c1);
DFFT DFFT_464__FPB_n1644(net1221,net585,net606_c1);
DFFT DFFT_456__FPB_n1636(net1220,net586,net607_c1);
DFFT DFFT_448__FPB_n1628(net1219,net587,net608_c1);
DFFT DFFT_392__FPB_n1572(net1218,net589,net618_c1);
DFFT DFFT_384__FPB_n1564(net1217,net590,net610_c1);
DFFT DFFT_376__FPB_n1556(net1216,net591,net611_c1);
DFFT DFFT_368__FPB_n1548(net1215,net108,net619_c1);
DFFT DFFT_296__FPB_n1476(net1214,net96,net614_c1);
DFFT DFFT_288__FPB_n1468(net1213,net595,net615_c1);
DFFT DFFT_537__FPB_n1717(net1630,net602,net620_c1);
DFFT DFFT_529__FPB_n1709(net1212,net603,net621_c1);
DFFT DFFT_481__FPB_n1661(net1211,net604,net634_c1);
DFFT DFFT_473__FPB_n1653(net1210,net605,net622_c1);
DFFT DFFT_465__FPB_n1645(net1209,net606,net623_c1);
DFFT DFFT_457__FPB_n1637(net1208,net2302,net624_c1);
DFFT DFFT_449__FPB_n1629(net1207,net608,net625_c1);
DFFT DFFT_393__FPB_n1573(net1206,net220,net635_c1);
DFFT DFFT_385__FPB_n1565(net1205,net2301,net636_c1);
DFFT DFFT_377__FPB_n1557(net1204,net611,net627_c1);
DFFT DFFT_369__FPB_n1549(net1203,net313,net628_c1);
DFFT DFFT_297__FPB_n1477(net1202,net614,net631_c1);
DFFT DFFT_289__FPB_n1469(net1201,net615,net632_c1);
DFFT DFFT_490__FPB_n1670(net1200,net715,net638_c1);
DFFT DFFT_482__FPB_n1662(net1199,net210,net639_c1);
DFFT DFFT_474__FPB_n1654(net1198,net622,net640_c1);
DFFT DFFT_466__FPB_n1646(net1197,net623,net641_c1);
DFFT DFFT_458__FPB_n1638(net1196,net624,net642_c1);
DFFT DFFT_394__FPB_n1574(net1195,net114,net645_c1);
DFFT DFFT_386__FPB_n1566(net1194,net230,net650_c1);
DFFT DFFT_378__FPB_n1558(net1193,net627,net646_c1);
DFFT DFFT_298__FPB_n1478(net1192,net2300,net651_c1);
XOR2T XOR2T_134_R0(net1958,net132,net665,net6_c1);
XOR2T XOR2T_44_n45(net1191,net51,net379,net46_c1);
XOR2T XOR2T_62_n63(net1190,net269,net288,net54_c1);
XOR2T XOR2T_47_n48(net2152,net256,net143,net62_c1);
XOR2T XOR2T_72_n73(net1189,net209,net392,net64_c1);
XOR2T XOR2T_65_n66(net1188,net76,net458,net71_c1);
XOR2T XOR2T_74_n75(net1187,net165,net177,net75_c1);
XOR2T XOR2T_91_n92(net1186,net195,net68,net78_c1);
XOR2T XOR2T_93_n94(net1185,net95,net559,net86_c1);
XOR2T XOR2T_89_n90(net1184,net73,net474,net68_c1);
AND2T AND2T_103_n104(net1183,net312,net391,net106_c1);
AND2T AND2T_112_n113(net1182,net105,net579,net107_c1);
AND2T AND2T_114_n115(net1181,net329,net600,net115_c1);
AND2T AND2T_106_n107(net1180,net121,net437,net116_c1);
AND2T AND2T_131_n132(net1179,net260,net472,net118_c1);
AND2T AND2T_123_n124(net1178,net150,net676,net119_c1);
AND2T AND2T_140_n141(net1177,net273,net634,net122_c1);
AND2T AND2T_132_n133(net1176,net232,net456,net123_c1);
AND2T AND2T_124_n125(net1175,net229,net705,net124_c1);
AND2T AND2T_116_n117(net1174,net129,net578,net125_c1);
AND2T AND2T_109_n110(net1173,net126,net557,net100_c1);
AND2T AND2T_141_n142(net1172,net207,net704,net127_c1);
AND2T AND2T_126_n127(net1171,net335,net390,net130_c1);
AND2T AND2T_118_n119(net1170,net226,net650,net131_c1);
AND2T AND2T_135_n136(net1959,net106,net675,net132_c1);
AND2T AND2T_129_n130(net1169,net222,net556,net109_c1);
DFFT DFFT_539__FPB_n1719(net1168,net157,net652_c1);
DFFT DFFT_491__FPB_n1671(net1167,net638,net653_c1);
DFFT DFFT_483__FPB_n1663(net1166,net639,net654_c1);
DFFT DFFT_475__FPB_n1655(net1165,net640,net655_c1);
DFFT DFFT_467__FPB_n1647(net1164,net641,net656_c1);
DFFT DFFT_459__FPB_n1639(net1163,net642,net665_c1);
DFFT DFFT_395__FPB_n1575(net1162,net645,net659_c1);
DFFT DFFT_387__FPB_n1567(net1161,net131,net660_c1);
DFFT DFFT_379__FPB_n1559(net1160,net646,net661_c1);
DFFT DFFT_299__FPB_n1479(net1159,net264,net663_c1);
DFFT DFFT_492__FPB_n1672(net1158,net653,net668_c1);
DFFT DFFT_484__FPB_n1664(net1157,net654,net669_c1);
DFFT DFFT_476__FPB_n1656(net1156,net655,net675_c1);
DFFT DFFT_468__FPB_n1648(net1155,net656,net670_c1);
DFFT DFFT_396__FPB_n1576(net1154,net659,net676_c1);
DFFT DFFT_388__FPB_n1568(net1153,net2299,net673_c1);
DFFT DFFT_511_Q3(net1152,net689,net9_c1);
DFFT DFFT_540_Q0(net1151,net652,net4_c1);
DFFT DFFT_527_Q2(net1150,net564,net7_c1);
DFFT DFFT_538_Q1(net1760,net620,net5_c1);
DFFT DFFT_493__FPB_n1673(net1149,net668,net679_c1);
DFFT DFFT_485__FPB_n1665(net1148,net669,net680_c1);
DFFT DFFT_477__FPB_n1657(net1147,net265,net681_c1);
DFFT DFFT_469__FPB_n1649(net2022,net670,net682_c1);
DFFT DFFT_397__FPB_n1577(net1146,net334,net685_c1);
DFFT DFFT_389__FPB_n1569(net1145,net673,net686_c1);
DFFT DFFT_494__FPB_n1674(net1144,net679,net691_c1);
DFFT DFFT_486__FPB_n1666(net1143,net680,net692_c1);
DFFT DFFT_478__FPB_n1658(net1142,net681,net693_c1);
DFFT DFFT_398__FPB_n1578(net1141,net2298,net695_c1);
DFFT DFFT_495__FPB_n1675(net1140,net691,net704_c1);
DFFT DFFT_487__FPB_n1667(net1139,net692,net699_c1);
DFFT DFFT_479__FPB_n1659(net1138,net693,net700_c1);
DFFT DFFT_399__FPB_n1579(net1137,net695,net705_c1);
AND2T AND2T_120_R3(net1136,net104,net110,net11_c1);
AND2T AND2T_23_n23(net1135,net19,net394,net21_c1);
AND2T AND2T_24_n24(net1134,net21,net408,net24_c1);
AND2T AND2T_33_n34(net1133,net180,net341,net31_c1);
AND2T AND2T_50_n51(net1132,net29,net56,net34_c1);
AND2T AND2T_42_n43(net1131,net30,net187,net35_c1);
AND2T AND2T_27_n27(net1130,net32,net285,net37_c1);
AND2T AND2T_19_n19(net1129,net339,net271,net38_c1);
AND2T AND2T_43_n44(net1128,net35,net25,net41_c1);
AND2T AND2T_35_n36(net1127,net47,net380,net42_c1);
AND2T AND2T_28_n28(net1126,net253,net2303,net43_c1);
AND2T AND2T_29_n30(net1125,net20,net350,net18_c1);
AND2T AND2T_61_n62(net1124,net153,net459,net49_c1);
AND2T AND2T_53_n54(net1123,net280,net477,net50_c1);
AND2T AND2T_54_n55(net1122,net238,net498,net55_c1);
AND2T AND2T_38_n39(net1121,net298,net406,net57_c1);
AND2T AND2T_49_n50(net1120,net67,net393,net29_c1);
AND2T AND2T_57_n58(net1119,net152,net281,net72_c1);
AND2T AND2T_82_n83(net1118,net79,net438,net74_c1);
AND2T AND2T_66_n67(net1117,net300,net198,net76_c1);
AND2T AND2T_59_n60(net1116,net44,net562,net39_c1);
AND2T AND2T_75_n76(net1115,net272,net422,net80_c1);
AND2T AND2T_67_n68(net1114,net242,net476,net81_c1);
AND2T AND2T_92_n93(net1113,net86,net293,net82_c1);
AND2T AND2T_76_n77(net1112,net178,net371,net84_c1);
AND2T AND2T_69_n70(net1111,net53,net582,net48_c1);
AND2T AND2T_85_n86(net1110,net83,net475,net87_c1);
AND2T AND2T_78_n79(net1109,net88,net327,net91_c1);
AND2T AND2T_95_n96(net1108,net328,net558,net92_c1);
AND2T AND2T_87_n88(net1107,net90,net541,net93_c1);
AND2T AND2T_88_n89(net1106,net204,net560,net95_c1);
DFFT DFFT_200__FPB_n1380(net1105,net599,net458_c1);
DFFT DFFT_496__FPB_n1676(net1104,net24,net708_c1);
DFFT DFFT_488__FPB_n1668(net1103,net699,net709_c1);
DFFT DFFT_201__FPB_n1381(net1102,net71,net476_c1);
DFFT DFFT_497__FPB_n1677(net1101,net708,net714_c1);
DFFT DFFT_489__FPB_n1669(net1100,net709,net715_c1);
DFFT DFFT_210__FPB_n1390(net1099,net2295,net494_c1);
DFFT DFFT_202__FPB_n1382(net1098,net193,net495_c1);
DFFT DFFT_498__FPB_n1678(net1097,net714,net720_c1);
OR2T OR2T_133_R1(net1096,net123,net118,net8_c1);
OR2T OR2T_127_R2(net1095,net130,net119,net10_c1);
OR2T OR2T_22_n22(net1094,net336,net274,net19_c1);
OR2T OR2T_30_n31(net1093,net237,net282,net20_c1);
OR2T OR2T_31_n32(net1092,net159,net356,net23_c1);
OR2T OR2T_40_n41(net1091,net297,net440,net25_c1);
OR2T OR2T_25_n25(net1090,net233,net246,net27_c1);
OR2T OR2T_41_n42(net1089,net199,net290,net30_c1);
OR2T OR2T_26_n26(net1088,net326,net171,net32_c1);
OR2T OR2T_34_n35(net1087,net31,net23,net36_c1);
OR2T OR2T_51_n52(net1086,net34,net46,net40_c1);
OR2T OR2T_60_n61(net1085,net279,net439,net44_c1);
OR2T OR2T_52_n53(net1084,net40,net303,net45_c1);
OR2T OR2T_36_n37(net1083,net286,net407,net47_c1);
OR2T OR2T_45_n46(net1082,net266,net423,net51_c1);
OR2T OR2T_37_n38(net1081,net292,net362,net52_c1);
OR2T OR2T_46_n47(net1080,net259,net478,net56_c1);
OR2T OR2T_39_n40(net1079,net338,net424,net22_c1);
OR2T OR2T_71_n72(net1078,net310,net637,net59_c1);
OR2T OR2T_63_n64(net1077,net49,net520,net60_c1);
OR2T OR2T_80_n81(net1076,net17,net404,net63_c1);
OR2T OR2T_64_n65(net1075,net60,net39,net65_c1);
OR2T OR2T_48_n49(net1074,net186,net499,net67_c1);
OR2T OR2T_81_n82(net1073,net194,net421,net69_c1);
OR2T OR2T_73_n74(net1072,net245,net405,net70_c1);
OR2T OR2T_90_n91(net1071,net166,net540,net73_c1);
OR2T OR2T_84_n85(net1070,net324,net457,net83_c1);
OR2T OR2T_68_n69(net1069,net139,net561,net85_c1);
OR2T OR2T_86_n87(net1068,net87,net497,net90_c1);
OR2T OR2T_79_n80(net1892,net306,net378,net58_c1);
OR2T OR2T_96_n97(net1067,net308,net601,net94_c1);
OR2T OR2T_98_n99(net1066,net192,net651,net97_c1);
DFFT DFFT_211__FPB_n1391(net1065,net494,net516_c1);
DFFT DFFT_203__FPB_n1383(net1064,net495,net517_c1);
DFFT DFFT_499__FPB_n1679(net1063,net720,net724_c1);
DFFT DFFT_220__FPB_n1400(net1062,net664,net343_c1);
DFFT DFFT_300__FPB_n1480(net1061,net663,net533_c1);
DFFT DFFT_212__FPB_n1392(net1060,net516,net536_c1);
DFFT DFFT_204__FPB_n1384(net1059,net517,net537_c1);
DFFT DFFT_221__FPB_n1401(net1058,net343,net344_c1);
DFFT DFFT_301__FPB_n1481(net1057,net533,net552_c1);
DFFT DFFT_213__FPB_n1393(net1056,net536,net554_c1);
DFFT DFFT_205__FPB_n1385(net1055,net537,net561_c1);
NOTT NOTT_20_n20(net1054,net283,net16_c1);
NOTT NOTT_21_n21(net1053,net302,net17_c1);
NOTT NOTT_32_n33(net1052,net179,net26_c1);
NOTT NOTT_17_n17(net1051,net270,net28_c1);
NOTT NOTT_18_n18(net1050,net261,net33_c1);
NOTT NOTT_70_n71(net1049,net81,net53_c1);
NOTT NOTT_55_n56(net1048,net299,net61_c1);
NOTT NOTT_56_n57(net1047,net251,net66_c1);
NOTT NOTT_58_n59(net1046,net243,net77_c1);
NOTT NOTT_83_n84(net1045,net320,net79_c1);
NOTT NOTT_77_n78(net1044,net301,net88_c1);
NOTT NOTT_94_n95(net1043,net82,net89_c1);
NOTT NOTT_97_n98(net1042,net94,net96_c1);
DFFT DFFT_230__FPB_n1410(net1041,net401,net345_c1);
DFFT DFFT_222__FPB_n1402(net1040,net344,net346_c1);
DFFT DFFT_150__FPB_n1330(net1039,net197,net347_c1);
DFFT DFFT_310__FPB_n1490(net1038,net688,net581_c1);
DFFT DFFT_302__FPB_n1482(net1037,net552,net572_c1);
DFFT DFFT_214__FPB_n1394(net1370,net554,net576_c1);
DFFT DFFT_206__FPB_n1386(net1036,net85,net582_c1);
XOR2T XOR2T_100_n101(net1035,net92,net677,net99_c1);
OR2T OR2T_102_n103(net1034,net93,net581,net103_c1);
OR2T OR2T_111_n112(net1500,net213,net580,net105_c1);
OR2T OR2T_113_n114(net1033,net325,net321,net111_c1);
XOR2T XOR2T_105_n106(net1032,net314,net420,net112_c1);
OR2T OR2T_130_n131(net1031,net134,net419,net113_c1);
XOR2T XOR2T_122_n123(net1030,net225,net635,net114_c1);
OR2T OR2T_115_n116(net1029,net115,net619,net120_c1);
OR2T OR2T_108_n109(net1028,net316,net473,net126_c1);
OR2T OR2T_125_n126(net1027,net124,net697,net128_c1);
XOR2T XOR2T_117_n118(net1026,net332,net636,net129_c1);
OR2T OR2T_119_n120(net1025,net254,net618,net104_c1);
XOR2T XOR2T_128_n129(net1024,net221,net217,net134_c1);
DFFT DFFT_231__FPB_n1411(net1371,net345,net348_c1);
DFFT DFFT_223__FPB_n1403(net1023,net346,net349_c1);
DFFT DFFT_151__FPB_n1331(net1696,net172,net350_c1);
DFFT DFFT_311__FPB_n1491(net1022,net206,net593_c1);
DFFT DFFT_303__FPB_n1483(net1021,net572,net594_c1);
DFFT DFFT_215__FPB_n1395(net1020,net576,net597_c1);
DFFT DFFT_207__FPB_n1387(net1019,net211,net598_c1);
DFFT DFFT_320__FPB_n1500(net1018,net703,net351_c1);
DFFT DFFT_240__FPB_n1420(net1017,net433,net352_c1);
DFFT DFFT_232__FPB_n1412(net1016,net348,net353_c1);
DFFT DFFT_224__FPB_n1404(net1015,net349,net354_c1);
DFFT DFFT_160__FPB_n1340(net1014,net436,net355_c1);
DFFT DFFT_152__FPB_n1332(net1697,net173,net356_c1);
DFFT DFFT_400__FPB_n1580(net1013,net196,net609_c1);
DFFT DFFT_312__FPB_n1492(net1012,net593,net612_c1);
DFFT DFFT_304__FPB_n1484(net1011,net594,net613_c1);
DFFT DFFT_216__FPB_n1396(net1010,net2297,net616_c1);
DFFT DFFT_208__FPB_n1388(net1009,net598,net617_c1);
DFFT DFFT_321__FPB_n1501(net1008,net351,net357_c1);
DFFT DFFT_241__FPB_n1421(net1007,net352,net358_c1);
DFFT DFFT_233__FPB_n1413(net1006,net2296,net359_c1);
DFFT DFFT_225__FPB_n1405(net1005,net354,net360_c1);
DFFT DFFT_161__FPB_n1341(net1004,net355,net362_c1);
DFFT DFFT_153__FPB_n1333(net1003,net250,net361_c1);
DFFT DFFT_401__FPB_n1581(net1002,net609,net626_c1);
DFFT DFFT_313__FPB_n1493(net1001,net612,net629_c1);
DFFT DFFT_305__FPB_n1485(net1000,net613,net630_c1);
DFFT DFFT_217__FPB_n1397(net999,net616,net637_c1);
DFFT DFFT_209__FPB_n1389(net998,net617,net633_c1);
AND2T AND2T_99_n100(net997,net331,net666,net98_c1);
DFFT DFFT_330__FPB_n1510(net996,net466,net363_c1);
DFFT DFFT_322__FPB_n1502(net995,net357,net364_c1);
DFFT DFFT_250__FPB_n1430(net994,net469,net365_c1);
DFFT DFFT_242__FPB_n1422(net993,net358,net371_c1);
DFFT DFFT_234__FPB_n1414(net992,net359,net366_c1);
DFFT DFFT_226__FPB_n1406(net991,net360,net367_c1);
DFFT DFFT_170__FPB_n1350(net990,net471,net368_c1);
DFFT DFFT_162__FPB_n1342(net989,net22,net369_c1);
DFFT DFFT_154__FPB_n1334(net988,net361,net370_c1);
DFFT DFFT_410__FPB_n1590(net987,net717,net643_c1);
DFFT DFFT_402__FPB_n1582(net986,net626,net644_c1);
DFFT DFFT_314__FPB_n1494(net985,net629,net647_c1);
DFFT DFFT_306__FPB_n1486(net984,net630,net648_c1);
DFFT DFFT_218__FPB_n1398(net983,net268,net649_c1);
DFFT DFFT_331__FPB_n1511(net982,net2294,net372_c1);
DFFT DFFT_323__FPB_n1503(net981,net364,net373_c1);
DFFT DFFT_251__FPB_n1431(net980,net365,net378_c1);
DFFT DFFT_243__FPB_n1423(net979,net191,net374_c1);
DFFT DFFT_235__FPB_n1415(net978,net366,net375_c1);
DFFT DFFT_227__FPB_n1407(net977,net367,net376_c1);
DFFT DFFT_171__FPB_n1351(net976,net368,net379_c1);
DFFT DFFT_163__FPB_n1343(net975,net369,net377_c1);
DFFT DFFT_155__FPB_n1335(net974,net370,net380_c1);
DFFT DFFT_411__FPB_n1591(net973,net643,net657_c1);
DFFT DFFT_403__FPB_n1583(net972,net644,net658_c1);
DFFT DFFT_315__FPB_n1495(net971,net647,net662_c1);
DFFT DFFT_307__FPB_n1487(net970,net648,net666_c1);
DFFT DFFT_219__FPB_n1399(net969,net649,net664_c1);
DFFT DFFT_420__FPB_n1600(net968,net725,net390_c1);
DFFT DFFT_340__FPB_n1520(net967,net510,net381_c1);
DFFT DFFT_332__FPB_n1512(net966,net372,net382_c1);
DFFT DFFT_324__FPB_n1504(net965,net373,net391_c1);
DFFT DFFT_260__FPB_n1440(net964,net515,net383_c1);
DFFT DFFT_252__FPB_n1432(net963,net257,net384_c1);
DFFT DFFT_244__FPB_n1424(net962,net374,net385_c1);
DFFT DFFT_236__FPB_n1416(net1893,net375,net386_c1);
DFFT DFFT_228__FPB_n1408(net961,net376,net392_c1);
DFFT DFFT_180__FPB_n1360(net960,net519,net393_c1);
DFFT DFFT_172__FPB_n1352(net959,net342,net387_c1);
DFFT DFFT_164__FPB_n1344(net958,net377,net388_c1);
DFFT DFFT_156__FPB_n1336(net957,net235,net389_c1);
DFFT DFFT_148__FPB_n1328(net956,net223,net394_c1);
DFFT DFFT_500__FPB_n1680(net955,net724,net667_c1);
DFFT DFFT_412__FPB_n1592(net954,net657,net671_c1);
DFFT DFFT_404__FPB_n1584(net953,net2293,net672_c1);
DFFT DFFT_316__FPB_n1496(net952,net662,net674_c1);
DFFT DFFT_308__FPB_n1488(net951,net98,net677_c1);
DFFT DFFT_421__FPB_n1601(net950,net311,net395_c1);
DFFT DFFT_341__FPB_n1521(net949,net381,net396_c1);
DFFT DFFT_333__FPB_n1513(net948,net382,net397_c1);
DFFT DFFT_325__FPB_n1505(net947,net33,net398_c1);
DFFT DFFT_261__FPB_n1441(net946,net383,net399_c1);
DFFT DFFT_253__FPB_n1433(net945,net384,net404_c1);
DFFT DFFT_245__FPB_n1425(net944,net385,net400_c1);
DFFT DFFT_237__FPB_n1417(net943,net386,net405_c1);
DFFT DFFT_229__FPB_n1409(net942,net247,net401_c1);
DFFT DFFT_181__FPB_n1361(net941,net170,net402_c1);
DFFT DFFT_173__FPB_n1353(net940,net387,net403_c1);
DFFT DFFT_165__FPB_n1345(net939,net388,net406_c1);
DFFT DFFT_157__FPB_n1337(net938,net389,net407_c1);
DFFT DFFT_149__FPB_n1329(net937,net278,net408_c1);
DFFT DFFT_501__FPB_n1681(net936,net2292,net678_c1);
DFFT DFFT_413__FPB_n1593(net935,net671,net683_c1);
DFFT DFFT_405__FPB_n1585(net934,net672,net684_c1);
DFFT DFFT_317__FPB_n1497(net933,net674,net687_c1);
DFFT DFFT_309__FPB_n1489(net932,net101,net688_c1);
DFFT DFFT_430__FPB_n1610(net931,net109,net419_c1);
DFFT DFFT_422__FPB_n1602(net930,net395,net409_c1);
DFFT DFFT_350__FPB_n1530(net929,net551,net410_c1);
DFFT DFFT_342__FPB_n1522(net928,net396,net411_c1);
DFFT DFFT_334__FPB_n1514(net927,net397,net420_c1);
DFFT DFFT_326__FPB_n1506(net926,net398,net412_c1);
DFFT DFFT_270__FPB_n1450(net925,net2285,net413_c1);
DFFT DFFT_262__FPB_n1442(net924,net399,net421_c1);
DFFT DFFT_254__FPB_n1434(net923,net248,net414_c1);
DFFT DFFT_246__FPB_n1426(net922,net400,net415_c1);
DFFT DFFT_238__FPB_n1418(net921,net75,net422_c1);
DFFT DFFT_190__FPB_n1370(net920,net276,net416_c1);
DFFT DFFT_182__FPB_n1362(net919,net402,net417_c1);
DFFT DFFT_174__FPB_n1354(net918,net403,net423_c1);
DFFT DFFT_166__FPB_n1346(net917,net151,net424_c1);
DFFT DFFT_158__FPB_n1338(net916,net330,net418_c1);
DFFT DFFT_510__FPB_n1690(net915,net729,net689_c1);
DFFT DFFT_502__FPB_n1682(net914,net678,net690_c1);
DFFT DFFT_414__FPB_n1594(net913,net683,net697_c1);
DFFT DFFT_406__FPB_n1586(net912,net684,net694_c1);
DFFT DFFT_318__FPB_n1498(net911,net687,net696_c1);
DFFT DFFT_142__FPB_n143(net910,net138,net732_c1);
DFFT DFFT_143__FPB_n144(net2153,net142,net733_c1);
SPLITT Split_600_n1780(net231,net202_c1,net307_c1);
SPLITT Split_601_n1781(net103,net207_c1,net312_c1);
DFFT DFFT_431__FPB_n1611(net909,net113,net425_c1);
DFFT DFFT_423__FPB_n1603(net908,net409,net426_c1);
DFFT DFFT_351__FPB_n1531(net907,net410,net427_c1);
DFFT DFFT_343__FPB_n1523(net906,net2291,net437_c1);
DFFT DFFT_335__FPB_n1515(net905,net318,net428_c1);
DFFT DFFT_327__FPB_n1507(net904,net412,net429_c1);
DFFT DFFT_271__FPB_n1451(net903,net413,net430_c1);
DFFT DFFT_263__FPB_n1443(net902,net227,net438_c1);
DFFT DFFT_255__FPB_n1435(net901,net414,net431_c1);
DFFT DFFT_247__FPB_n1427(net900,net415,net432_c1);
DFFT DFFT_239__FPB_n1419(net899,net80,net433_c1);
DFFT DFFT_191__FPB_n1371(net898,net416,net439_c1);
DFFT DFFT_183__FPB_n1363(net897,net417,net434_c1);
DFFT DFFT_175__FPB_n1355(net896,net147,net435_c1);
DFFT DFFT_167__FPB_n1347(net895,net224,net440_c1);
DFFT DFFT_159__FPB_n1339(net894,net418,net436_c1);
DFFT DFFT_503__FPB_n1683(net893,net690,net698_c1);
DFFT DFFT_415__FPB_n1595(net892,net214,net701_c1);
DFFT DFFT_407__FPB_n1587(net891,net694,net702_c1);
DFFT DFFT_319__FPB_n1499(net890,net696,net703_c1);
SPLITT Split_602_n1782(net116,net213_c1,net316_c1);
SPLITT Split_610_n1790(net234,net211_c1,net317_c1);
SPLITT Split_603_n1783(net100,net217_c1,net321_c1);
SPLITT Split_611_n1791(net135,net215_c1,net322_c1);
SPLITT Split_620_n1800(net122,net137_c1,net240_c1);
SPLITT Split_604_n1784(net107,net221_c1,net325_c1);
SPLITT Split_612_n1792(net322,net223_c1,net326_c1);
SPLITT Split_541_n1721(net15,net138_c1,net241_c1);
SPLITT Split_621_n1801(net240,net139_c1,net242_c1);
DFFT DFFT_144__FPB_n145(net889,net175,net734_c1);
SPLITT Split_605_n1785(net111,net225_c1,net329_c1);
SPLITT Split_613_n1793(net215,net224_c1,net330_c1);
SPLITT Split_542_n1722(net14,net142_c1,net243_c1);
SPLITT Split_550_n1730(net284,net140_c1,net244_c1);
SPLITT Split_622_n1802(net137,net141_c1,net245_c1);
SPLITT Split_630_n1810(net289,net143_c1,net246_c1);
SPLITT Split_606_n1786(net120,net229_c1,net332_c1);
SPLITT Split_614_n1794(net136,net228_c1,net333_c1);
SPLITT Split_543_n1723(net13,net146_c1,net247_c1);
SPLITT Split_551_n1731(net182,net145_c1,net248_c1);
SPLITT Split_623_n1803(net127,net144_c1,net249_c1);
SPLITT Split_631_n1811(net181,net147_c1,net250_c1);
SPLITT Split_607_n1787(net128,net232_c1,net335_c1);
SPLITT Split_615_n1795(net333,net233_c1,net336_c1);
SPLITT Split_544_n1724(net146,net151_c1,net251_c1);
SPLITT Split_552_n1732(net0,net149_c1,net252_c1);
SPLITT Split_560_n1740(net37,net153_c1,net253_c1);
SPLITT Split_624_n1804(net249,net150_c1,net254_c1);
SPLITT Split_632_n1812(net734,net148_c1,net255_c1);
SPLITT Split_640_n1820(net188,net152_c1,net256_c1);
SPLITT Split_608_n1788(net133,net234_c1,net337_c1);
SPLITT Split_616_n1796(net228,net235_c1,net338_c1);
SPLITT Split_545_n1725(net12,net155_c1,net257_c1);
SPLITT Split_553_n1733(net149,net156_c1,net258_c1);
SPLITT Split_561_n1741(net43,net158_c1,net259_c1);
SPLITT Split_625_n1805(net144,net157_c1,net260_c1);
SPLITT Split_633_n1813(net255,net159_c1,net261_c1);
SPLITT Split_641_n1821(net737,net154_c1,net262_c1);
SPLITT Split_609_n1789(net337,net237_c1,net339_c1);
SPLITT Split_617_n1797(net117,net236_c1,net340_c1);
SPLITT Split_546_n1726(net3,net164_c1,net263_c1);
SPLITT Split_554_n1734(net28,net162_c1,net264_c1);
SPLITT Split_562_n1742(net18,net161_c1,net265_c1);
SPLITT Split_570_n1750(net208,net166_c1,net266_c1);
SPLITT Split_626_n1806(net732,net160_c1,net267_c1);
SPLITT Split_634_n1814(net148,net163_c1,net268_c1);
SPLITT Split_642_n1822(net262,net165_c1,net269_c1);
SPLITT Split_618_n1798(net340,net238_c1,net341_c1);
SPLITT Split_547_n1727(net164,net173_c1,net270_c1);
SPLITT Split_555_n1735(net162,net172_c1,net271_c1);
SPLITT Split_563_n1743(net161,net170_c1,net272_c1);
SPLITT Split_571_n1751(net45,net169_c1,net273_c1);
SPLITT Split_627_n1807(net267,net171_c1,net274_c1);
SPLITT Split_635_n1815(net735,net167_c1,net275_c1);
SPLITT Split_643_n1823(net154,net168_c1,net276_c1);
SPLITT Split_619_n1799(net236,net239_c1,net342_c1);
SPLITT Split_548_n1728(net2,net175_c1,net277_c1);
SPLITT Split_556_n1736(net38,net174_c1,net278_c1);
SPLITT Split_564_n1744(net36,net176_c1,net279_c1);
SPLITT Split_572_n1752(net169,net178_c1,net280_c1);
SPLITT Split_580_n1760(net216,net177_c1,net281_c1);
SPLITT Split_628_n1808(net160,net179_c1,net282_c1);
SPLITT Split_636_n1816(net275,net180_c1,net283_c1);
SPLITT Split_549_n1729(net1,net182_c1,net284_c1);
SPLITT Split_557_n1737(net174,net187_c1,net285_c1);
SPLITT Split_565_n1745(net176,net186_c1,net286_c1);
SPLITT Split_573_n1753(net50,net183_c1,net287_c1);
SPLITT Split_581_n1761(net77,net184_c1,net288_c1);
SPLITT Split_629_n1809(net733,net181_c1,net289_c1);
SPLITT Split_637_n1817(net167,net185_c1,net290_c1);
SPLITT Split_558_n1738(net16,net191_c1,net291_c1);
SPLITT Split_566_n1746(net42,net193_c1,net292_c1);
SPLITT Split_574_n1754(net183,net192_c1,net293_c1);
SPLITT Split_582_n1762(net65,net190_c1,net294_c1);
SPLITT Split_590_n1770(net84,net189_c1,net295_c1);
SPLITT Split_638_n1818(net736,net188_c1,net296_c1);
SPLITT Split_559_n1739(net27,net197_c1,net297_c1);
SPLITT Split_567_n1747(net52,net198_c1,net298_c1);
SPLITT Split_575_n1755(net55,net196_c1,net299_c1);
SPLITT Split_583_n1763(net190,net195_c1,net300_c1);
SPLITT Split_591_n1771(net189,net194_c1,net301_c1);
SPLITT Split_639_n1819(net296,net199_c1,net302_c1);
SPLITT Split_568_n1748(net57,net204_c1,net303_c1);
SPLITT Split_576_n1756(net61,net201_c1,net304_c1);
SPLITT Split_584_n1764(net48,net200_c1,net305_c1);
SPLITT Split_592_n1772(net91,net203_c1,net306_c1);
SPLITT Split_569_n1749(net41,net208_c1,net308_c1);
SPLITT Split_577_n1757(net304,net206_c1,net309_c1);
SPLITT Split_585_n1765(net305,net209_c1,net310_c1);
SPLITT Split_593_n1773(net63,net205_c1,net311_c1);
SPLITT Split_578_n1758(net201,net210_c1,net313_c1);
SPLITT Split_586_n1766(net200,net214_c1,net314_c1);
SPLITT Split_594_n1774(net205,net212_c1,net315_c1);
SPLITT Split_579_n1759(net66,net216_c1,net318_c1);
SPLITT Split_587_n1767(net59,net218_c1,net319_c1);
SPLITT Split_595_n1775(net69,net219_c1,net320_c1);
SPLITT Split_588_n1768(net64,net220_c1,net323_c1);
SPLITT Split_596_n1776(net74,net222_c1,net324_c1);
DFFT DFFT_145__FPB_n146(net888,net140,net735_c1);
SPLITT Split_589_n1769(net70,net227_c1,net327_c1);
SPLITT Split_597_n1777(net89,net226_c1,net328_c1);
SPLITT Split_598_n1778(net97,net230_c1,net331_c1);
SPLITT Split_599_n1779(net99,net231_c1,net334_c1);
DFFT DFFT_520__FPB_n1700(net887,net731,net441_c1);
DFFT DFFT_440__FPB_n1620(net886,net588,net456_c1);
DFFT DFFT_432__FPB_n1612(net885,net425,net442_c1);
DFFT DFFT_424__FPB_n1604(net884,net426,net443_c1);
DFFT DFFT_360__FPB_n1540(net883,net592,net444_c1);
DFFT DFFT_352__FPB_n1532(net882,net427,net445_c1);
DFFT DFFT_344__FPB_n1524(net881,net295,net446_c1);
DFFT DFFT_336__FPB_n1516(net880,net428,net447_c1);
DFFT DFFT_328__FPB_n1508(net879,net429,net448_c1);
DFFT DFFT_280__FPB_n1460(net878,net596,net449_c1);
DFFT DFFT_272__FPB_n1452(net877,net430,net457_c1);
DFFT DFFT_264__FPB_n1444(net876,net212,net450_c1);
DFFT DFFT_256__FPB_n1436(net875,net431,net451_c1);
DFFT DFFT_248__FPB_n1428(net874,net432,net452_c1);
DFFT DFFT_192__FPB_n1372(net1761,net54,net459_c1);
DFFT DFFT_184__FPB_n1364(net873,net434,net453_c1);
DFFT DFFT_176__FPB_n1356(net872,net435,net454_c1);
DFFT DFFT_168__FPB_n1348(net871,net317,net455_c1);
DFFT DFFT_512__FPB_n1692(net870,net158,net706_c1);
DFFT DFFT_504__FPB_n1684(net869,net698,net707_c1);
DFFT DFFT_416__FPB_n1596(net868,net701,net710_c1);
DFFT DFFT_408__FPB_n1588(net867,net702,net711_c1);
DFFT DFFT_146__FPB_n147(net866,net156,net736_c1);
DFFT DFFT_147__FPB_n148(net865,net252,net737_c1);
DFFT DFFT_521__FPB_n1701(net864,net441,net460_c1);
DFFT DFFT_441__FPB_n1621(net863,net155,net461_c1);
DFFT DFFT_433__FPB_n1613(net862,net442,net472_c1);
DFFT DFFT_425__FPB_n1605(net861,net443,net462_c1);
DFFT DFFT_361__FPB_n1541(net860,net444,net463_c1);
DFFT DFFT_353__FPB_n1533(net1501,net445,net464_c1);
DFFT DFFT_345__FPB_n1525(net859,net446,net473_c1);
DFFT DFFT_337__FPB_n1517(net858,net447,net465_c1);
DFFT DFFT_329__FPB_n1509(net857,net448,net466_c1);
DFFT DFFT_281__FPB_n1461(net856,net449,net474_c1);
DFFT DFFT_273__FPB_n1453(net855,net58,net475_c1);
DFFT DFFT_265__FPB_n1445(net854,net450,net467_c1);
DFFT DFFT_257__FPB_n1437(net853,net451,net468_c1);
DFFT DFFT_249__FPB_n1429(net852,net452,net469_c1);
DFFT DFFT_193__FPB_n1373(net851,net185,net470_c1);
DFFT DFFT_185__FPB_n1365(net850,net453,net477_c1);
DFFT DFFT_177__FPB_n1357(net849,net2290,net478_c1);
DFFT DFFT_169__FPB_n1349(net848,net455,net471_c1);
DFFT DFFT_513__FPB_n1693(net847,net706,net712_c1);
DFFT DFFT_505__FPB_n1685(net846,net707,net713_c1);
DFFT DFFT_417__FPB_n1597(net845,net710,net716_c1);
DFFT DFFT_409__FPB_n1589(net844,net711,net717_c1);
DFFT DFFT_530__FPB_n1710(net843,net621,net479_c1);
DFFT DFFT_522__FPB_n1702(net1631,net460,net480_c1);
DFFT DFFT_450__FPB_n1630(net842,net625,net481_c1);
DFFT DFFT_442__FPB_n1622(net841,net461,net482_c1);
DFFT DFFT_434__FPB_n1614(net840,net203,net483_c1);
DFFT DFFT_426__FPB_n1606(net839,net462,net484_c1);
DFFT DFFT_370__FPB_n1550(net838,net628,net485_c1);
DFFT DFFT_362__FPB_n1542(net837,net463,net486_c1);
DFFT DFFT_354__FPB_n1534(net836,net464,net487_c1);
DFFT DFFT_346__FPB_n1526(net835,net145,net488_c1);
DFFT DFFT_338__FPB_n1518(net834,net465,net489_c1);
DFFT DFFT_290__FPB_n1470(net833,net632,net490_c1);
DFFT DFFT_282__FPB_n1462(net832,net239,net491_c1);
DFFT DFFT_274__FPB_n1454(net831,net323,net497_c1);
DFFT DFFT_266__FPB_n1446(net830,net467,net492_c1);
DFFT DFFT_258__FPB_n1438(net829,net468,net493_c1);
DFFT DFFT_194__FPB_n1374(net828,net470,net496_c1);
DFFT DFFT_186__FPB_n1366(net827,net263,net498_c1);
DFFT DFFT_178__FPB_n1358(net826,net62,net499_c1);
DFFT DFFT_514__FPB_n1694(net825,net2289,net718_c1);
DFFT DFFT_506__FPB_n1686(net824,net713,net719_c1);
DFFT DFFT_418__FPB_n1598(net823,net716,net721_c1);
NOTT NOTT_101_n102(net822,net307,net101_c1);
NOTT NOTT_110_n111(net821,net315,net102_c1);
NOTT NOTT_104_n105(net820,net319,net108_c1);
NOTT NOTT_121_n122(net1437,net125,net110_c1);
NOTT NOTT_107_n108(net819,net287,net121_c1);
NOTT NOTT_136_n137(net818,net277,net133_c1);
NOTT NOTT_137_n138(net817,net244,net135_c1);
NOTT NOTT_138_n139(net816,net258,net136_c1);
NOTT NOTT_139_n140(net815,net241,net117_c1);
DFFT DFFT_531__FPB_n1711(net814,net479,net500_c1);
DFFT DFFT_523__FPB_n1703(net813,net480,net501_c1);
DFFT DFFT_451__FPB_n1631(net812,net481,net502_c1);
DFFT DFFT_443__FPB_n1623(net811,net482,net503_c1);
DFFT DFFT_435__FPB_n1615(net810,net483,net504_c1);
DFFT DFFT_427__FPB_n1607(net809,net2288,net505_c1);
DFFT DFFT_371__FPB_n1551(net808,net485,net506_c1);
DFFT DFFT_363__FPB_n1543(net807,net486,net507_c1);
DFFT DFFT_355__FPB_n1535(net806,net487,net508_c1);
DFFT DFFT_347__FPB_n1527(net805,net488,net509_c1);
DFFT DFFT_339__FPB_n1519(net804,net489,net510_c1);
DFFT DFFT_291__FPB_n1471(net803,net2287,net511_c1);
DFFT DFFT_283__FPB_n1463(net802,net491,net512_c1);
DFFT DFFT_275__FPB_n1455(net801,net218,net513_c1);
DFFT DFFT_267__FPB_n1447(net800,net492,net514_c1);
DFFT DFFT_259__FPB_n1439(net799,net493,net515_c1);
DFFT DFFT_195__FPB_n1375(net798,net2286,net520_c1);
DFFT DFFT_187__FPB_n1367(net797,net184,net518_c1);
DFFT DFFT_179__FPB_n1359(net796,net291,net519_c1);
DFFT DFFT_515__FPB_n1695(net795,net718,net722_c1);
DFFT DFFT_507__FPB_n1687(net794,net719,net723_c1);
DFFT DFFT_419__FPB_n1599(net793,net721,net725_c1);
DFFT DFFT_532__FPB_n1712(net792,net500,net521_c1);
DFFT DFFT_524__FPB_n1704(net791,net501,net522_c1);
DFFT DFFT_460__FPB_n1640(net790,net168,net523_c1);
DFFT DFFT_452__FPB_n1632(net789,net502,net524_c1);
DFFT DFFT_444__FPB_n1624(net788,net503,net525_c1);
DFFT DFFT_436__FPB_n1616(net787,net504,net526_c1);
DFFT DFFT_428__FPB_n1608(net786,net505,net527_c1);
DFFT DFFT_380__FPB_n1560(net785,net661,net528_c1);
DFFT DFFT_372__FPB_n1552(net784,net506,net529_c1);
DFFT DFFT_364__FPB_n1544(net783,net507,net530_c1);
DFFT DFFT_356__FPB_n1536(net782,net508,net531_c1);
DFFT DFFT_348__FPB_n1528(net781,net509,net532_c1);
DFFT DFFT_292__FPB_n1472(net780,net511,net534_c1);
DFFT DFFT_284__FPB_n1464(net779,net512,net540_c1);
DFFT DFFT_276__FPB_n1456(net778,net513,net541_c1);
DFFT DFFT_268__FPB_n1448(net777,net514,net535_c1);
DFFT DFFT_196__FPB_n1376(net776,net72,net538_c1);
DFFT DFFT_188__FPB_n1368(net2282,net518,net539_c1);
DFFT DFFT_516__FPB_n1696(net775,net722,net726_c1);
DFFT DFFT_508__FPB_n1688(net774,net723,net727_c1);
DFFT DFFT_533__FPB_n1713(net773,net521,net542_c1);
DFFT DFFT_525__FPB_n1705(net772,net522,net543_c1);
DFFT DFFT_461__FPB_n1641(net2219,net523,net544_c1);
DFFT DFFT_453__FPB_n1633(net771,net524,net545_c1);
DFFT DFFT_445__FPB_n1625(net770,net525,net546_c1);
DFFT DFFT_437__FPB_n1617(net769,net526,net547_c1);
DFFT DFFT_429__FPB_n1609(net768,net527,net556_c1);
DFFT DFFT_381__FPB_n1561(net767,net528,net548_c1);
DFFT DFFT_373__FPB_n1553(net766,net529,net549_c1);
DFFT DFFT_365__FPB_n1545(net765,net530,net550_c1);
DFFT DFFT_357__FPB_n1537(net764,net531,net557_c1);
DFFT DFFT_349__FPB_n1529(net763,net532,net551_c1);
DFFT DFFT_293__FPB_n1473(net762,net534,net558_c1);
DFFT DFFT_285__FPB_n1465(net761,net78,net559_c1);
DFFT DFFT_277__FPB_n1457(net760,net294,net560_c1);
DFFT DFFT_269__FPB_n1449(net759,net535,net553_c1);
DFFT DFFT_197__FPB_n1377(net758,net538,net555_c1);
DFFT DFFT_189__FPB_n1369(net2283,net539,net562_c1);
DFFT DFFT_517__FPB_n1697(net757,net726,net728_c1);
DFFT DFFT_509__FPB_n1689(net756,net727,net729_c1);
DFFT DFFT_534__FPB_n1714(net755,net542,net563_c1);
DFFT DFFT_526__FPB_n1706(net754,net543,net564_c1);
DFFT DFFT_470__FPB_n1650(net2023,net682,net565_c1);
DFFT DFFT_462__FPB_n1642(net753,net544,net566_c1);
DFFT DFFT_454__FPB_n1634(net752,net545,net567_c1);
DFFT DFFT_446__FPB_n1626(net751,net546,net568_c1);
DFFT DFFT_438__FPB_n1618(net750,net547,net569_c1);
DFFT DFFT_390__FPB_n1570(net749,net686,net570_c1);
DFFT DFFT_382__FPB_n1562(net748,net548,net578_c1);
DFFT DFFT_374__FPB_n1554(net747,net549,net571_c1);
DFFT DFFT_366__FPB_n1546(net746,net550,net579_c1);
DFFT DFFT_358__FPB_n1538(net745,net219,net580_c1);
DFFT DFFT_294__FPB_n1474(net744,net26,net573_c1);
DFFT DFFT_286__FPB_n1466(net743,net309,net574_c1);
DFFT DFFT_278__FPB_n1458(net742,net163,net575_c1);
DFFT DFFT_198__FPB_n1378(net741,net555,net577_c1);
DFFT DFFT_518__FPB_n1698(net740,net728,net730_c1);
SPLITT SplitCLK_4_525(net2281,net2282_c1,net2283_c1);
SPLITT SplitCLK_6_526(net2276,net2281_c1,net2280_c1);
SPLITT SplitCLK_2_527(net2277,net2279_c1,net2278_c1);
SPLITT SplitCLK_4_528(net2268,net2277_c1,net2276_c1);
SPLITT SplitCLK_6_529(net2270,net2275_c1,net2274_c1);
SPLITT SplitCLK_4_530(net2271,net2272_c1,net2273_c1);
SPLITT SplitCLK_2_531(net2269,net2270_c1,net2271_c1);
SPLITT SplitCLK_6_532(net2252,net2268_c1,net2269_c1);
SPLITT SplitCLK_0_533(net2262,net2267_c1,net2266_c1);
SPLITT SplitCLK_6_534(net2263,net2264_c1,net2265_c1);
SPLITT SplitCLK_4_535(net2254,net2263_c1,net2262_c1);
SPLITT SplitCLK_4_536(net2256,net2261_c1,net2260_c1);
SPLITT SplitCLK_2_537(net2257,net2258_c1,net2259_c1);
SPLITT SplitCLK_6_538(net2255,net2256_c1,net2257_c1);
SPLITT SplitCLK_4_539(net2253,net2255_c1,net2254_c1);
SPLITT SplitCLK_0_540(net2220,net2252_c1,net2253_c1);
SPLITT SplitCLK_6_541(net2246,net2250_c1,net2251_c1);
SPLITT SplitCLK_4_542(net2247,net2249_c1,net2248_c1);
SPLITT SplitCLK_4_543(net2238,net2246_c1,net2247_c1);
SPLITT SplitCLK_6_544(net2240,net2245_c1,net2244_c1);
SPLITT SplitCLK_6_545(net2241,net2242_c1,net2243_c1);
SPLITT SplitCLK_6_546(net2239,net2240_c1,net2241_c1);
SPLITT SplitCLK_6_547(net2222,net2238_c1,net2239_c1);
SPLITT SplitCLK_6_548(net2232,net2237_c1,net2236_c1);
SPLITT SplitCLK_4_549(net2233,net2234_c1,net2235_c1);
SPLITT SplitCLK_4_550(net2224,net2232_c1,net2233_c1);
SPLITT SplitCLK_6_551(net2226,net2230_c1,net2231_c1);
SPLITT SplitCLK_4_552(net2227,net2228_c1,net2229_c1);
SPLITT SplitCLK_6_553(net2225,net2227_c1,net2226_c1);
SPLITT SplitCLK_4_554(net2223,net2225_c1,net2224_c1);
SPLITT SplitCLK_2_555(net2221,net2223_c1,net2222_c1);
SPLITT SplitCLK_6_556(net2154,net2220_c1,net2221_c1);
SPLITT SplitCLK_4_557(net2217,net2219_c1,net2218_c1);
SPLITT SplitCLK_0_558(net2212,net2216_c1,net2217_c1);
SPLITT SplitCLK_6_559(net2213,net2215_c1,net2214_c1);
SPLITT SplitCLK_4_560(net2204,net2213_c1,net2212_c1);
SPLITT SplitCLK_6_561(net2206,net2210_c1,net2211_c1);
SPLITT SplitCLK_2_562(net2207,net2209_c1,net2208_c1);
SPLITT SplitCLK_6_563(net2205,net2206_c1,net2207_c1);
SPLITT SplitCLK_6_564(net2188,net2204_c1,net2205_c1);
SPLITT SplitCLK_4_565(net2198,net2202_c1,net2203_c1);
SPLITT SplitCLK_4_566(net2199,net2200_c1,net2201_c1);
SPLITT SplitCLK_0_567(net2190,net2198_c1,net2199_c1);
SPLITT SplitCLK_4_568(net2192,net2196_c1,net2197_c1);
SPLITT SplitCLK_4_569(net2193,net2195_c1,net2194_c1);
SPLITT SplitCLK_2_570(net2191,net2192_c1,net2193_c1);
SPLITT SplitCLK_0_571(net2189,net2190_c1,net2191_c1);
SPLITT SplitCLK_4_572(net2156,net2189_c1,net2188_c1);
SPLITT SplitCLK_6_573(net2182,net2187_c1,net2186_c1);
SPLITT SplitCLK_4_574(net2183,net2184_c1,net2185_c1);
SPLITT SplitCLK_4_575(net2174,net2182_c1,net2183_c1);
SPLITT SplitCLK_6_576(net2176,net2181_c1,net2180_c1);
SPLITT SplitCLK_4_577(net2177,net2179_c1,net2178_c1);
SPLITT SplitCLK_2_578(net2175,net2177_c1,net2176_c1);
SPLITT SplitCLK_2_579(net2158,net2174_c1,net2175_c1);
SPLITT SplitCLK_6_580(net2168,net2173_c1,net2172_c1);
SPLITT SplitCLK_4_581(net2169,net2171_c1,net2170_c1);
SPLITT SplitCLK_0_582(net2160,net2168_c1,net2169_c1);
SPLITT SplitCLK_6_583(net2162,net2167_c1,net2166_c1);
SPLITT SplitCLK_4_584(net2163,net2164_c1,net2165_c1);
SPLITT SplitCLK_2_585(net2161,net2163_c1,net2162_c1);
SPLITT SplitCLK_4_586(net2159,net2161_c1,net2160_c1);
SPLITT SplitCLK_2_587(net2157,net2159_c1,net2158_c1);
SPLITT SplitCLK_4_588(net2155,net2157_c1,net2156_c1);
SPLITT SplitCLK_0_589(net2024,net2154_c1,net2155_c1);
SPLITT SplitCLK_4_590(net2151,net2152_c1,net2153_c1);
SPLITT SplitCLK_6_591(net2146,net2151_c1,net2150_c1);
SPLITT SplitCLK_4_592(net2147,net2149_c1,net2148_c1);
SPLITT SplitCLK_0_593(net2138,net2146_c1,net2147_c1);
SPLITT SplitCLK_6_594(net2140,net2144_c1,net2145_c1);
SPLITT SplitCLK_4_595(net2141,net2142_c1,net2143_c1);
SPLITT SplitCLK_6_596(net2139,net2141_c1,net2140_c1);
SPLITT SplitCLK_6_597(net2122,net2138_c1,net2139_c1);
SPLITT SplitCLK_4_598(net2132,net2136_c1,net2137_c1);
SPLITT SplitCLK_4_599(net2133,net2135_c1,net2134_c1);
SPLITT SplitCLK_0_600(net2124,net2132_c1,net2133_c1);
SPLITT SplitCLK_6_601(net2126,net2131_c1,net2130_c1);
SPLITT SplitCLK_6_602(net2127,net2128_c1,net2129_c1);
SPLITT SplitCLK_4_603(net2125,net2127_c1,net2126_c1);
SPLITT SplitCLK_4_604(net2123,net2125_c1,net2124_c1);
SPLITT SplitCLK_0_605(net2090,net2122_c1,net2123_c1);
SPLITT SplitCLK_6_606(net2116,net2121_c1,net2120_c1);
SPLITT SplitCLK_0_607(net2117,net2118_c1,net2119_c1);
SPLITT SplitCLK_0_608(net2108,net2116_c1,net2117_c1);
SPLITT SplitCLK_6_609(net2110,net2115_c1,net2114_c1);
SPLITT SplitCLK_4_610(net2111,net2113_c1,net2112_c1);
SPLITT SplitCLK_6_611(net2109,net2111_c1,net2110_c1);
SPLITT SplitCLK_6_612(net2092,net2108_c1,net2109_c1);
SPLITT SplitCLK_2_613(net2102,net2106_c1,net2107_c1);
SPLITT SplitCLK_4_614(net2103,net2105_c1,net2104_c1);
SPLITT SplitCLK_4_615(net2094,net2102_c1,net2103_c1);
SPLITT SplitCLK_6_616(net2096,net2100_c1,net2101_c1);
SPLITT SplitCLK_4_617(net2097,net2098_c1,net2099_c1);
SPLITT SplitCLK_6_618(net2095,net2097_c1,net2096_c1);
SPLITT SplitCLK_4_619(net2093,net2095_c1,net2094_c1);
SPLITT SplitCLK_6_620(net2091,net2093_c1,net2092_c1);
SPLITT SplitCLK_6_621(net2026,net2090_c1,net2091_c1);
SPLITT SplitCLK_0_622(net2084,net2089_c1,net2088_c1);
SPLITT SplitCLK_4_623(net2085,net2086_c1,net2087_c1);
SPLITT SplitCLK_4_624(net2076,net2084_c1,net2085_c1);
SPLITT SplitCLK_6_625(net2078,net2082_c1,net2083_c1);
SPLITT SplitCLK_4_626(net2079,net2080_c1,net2081_c1);
SPLITT SplitCLK_6_627(net2077,net2079_c1,net2078_c1);
SPLITT SplitCLK_6_628(net2060,net2076_c1,net2077_c1);
SPLITT SplitCLK_0_629(net2070,net2074_c1,net2075_c1);
SPLITT SplitCLK_4_630(net2071,net2073_c1,net2072_c1);
SPLITT SplitCLK_4_631(net2062,net2071_c1,net2070_c1);
SPLITT SplitCLK_0_632(net2064,net2068_c1,net2069_c1);
SPLITT SplitCLK_4_633(net2065,net2067_c1,net2066_c1);
SPLITT SplitCLK_2_634(net2063,net2065_c1,net2064_c1);
SPLITT SplitCLK_4_635(net2061,net2063_c1,net2062_c1);
SPLITT SplitCLK_0_636(net2028,net2060_c1,net2061_c1);
SPLITT SplitCLK_6_637(net2054,net2058_c1,net2059_c1);
SPLITT SplitCLK_2_638(net2055,net2056_c1,net2057_c1);
SPLITT SplitCLK_4_639(net2046,net2055_c1,net2054_c1);
SPLITT SplitCLK_4_640(net2048,net2053_c1,net2052_c1);
SPLITT SplitCLK_4_641(net2049,net2051_c1,net2050_c1);
SPLITT SplitCLK_6_642(net2047,net2048_c1,net2049_c1);
SPLITT SplitCLK_6_643(net2030,net2046_c1,net2047_c1);
SPLITT SplitCLK_4_644(net2040,net2045_c1,net2044_c1);
SPLITT SplitCLK_4_645(net2041,net2043_c1,net2042_c1);
SPLITT SplitCLK_0_646(net2032,net2040_c1,net2041_c1);
SPLITT SplitCLK_6_647(net2034,net2039_c1,net2038_c1);
SPLITT SplitCLK_6_648(net2035,net2037_c1,net2036_c1);
SPLITT SplitCLK_4_649(net2033,net2035_c1,net2034_c1);
SPLITT SplitCLK_4_650(net2031,net2033_c1,net2032_c1);
SPLITT SplitCLK_2_651(net2029,net2031_c1,net2030_c1);
SPLITT SplitCLK_4_652(net2027,net2029_c1,net2028_c1);
SPLITT SplitCLK_2_653(net2025,net2027_c1,net2026_c1);
SPLITT SplitCLK_6_654(net1762,net2024_c1,net2025_c1);
SPLITT SplitCLK_4_655(net2021,net2023_c1,net2022_c1);
SPLITT SplitCLK_6_656(net2016,net2021_c1,net2020_c1);
SPLITT SplitCLK_4_657(net2017,net2018_c1,net2019_c1);
SPLITT SplitCLK_0_658(net2008,net2016_c1,net2017_c1);
SPLITT SplitCLK_0_659(net2010,net2015_c1,net2014_c1);
SPLITT SplitCLK_6_660(net2011,net2012_c1,net2013_c1);
SPLITT SplitCLK_2_661(net2009,net2010_c1,net2011_c1);
SPLITT SplitCLK_6_662(net1992,net2008_c1,net2009_c1);
SPLITT SplitCLK_0_663(net2002,net2007_c1,net2006_c1);
SPLITT SplitCLK_4_664(net2003,net2005_c1,net2004_c1);
SPLITT SplitCLK_4_665(net1994,net2002_c1,net2003_c1);
SPLITT SplitCLK_0_666(net1996,net2000_c1,net2001_c1);
SPLITT SplitCLK_0_667(net1997,net1999_c1,net1998_c1);
SPLITT SplitCLK_6_668(net1995,net1996_c1,net1997_c1);
SPLITT SplitCLK_4_669(net1993,net1995_c1,net1994_c1);
SPLITT SplitCLK_0_670(net1960,net1992_c1,net1993_c1);
SPLITT SplitCLK_0_671(net1986,net1990_c1,net1991_c1);
SPLITT SplitCLK_4_672(net1987,net1989_c1,net1988_c1);
SPLITT SplitCLK_4_673(net1978,net1986_c1,net1987_c1);
SPLITT SplitCLK_6_674(net1980,net1984_c1,net1985_c1);
SPLITT SplitCLK_4_675(net1981,net1983_c1,net1982_c1);
SPLITT SplitCLK_6_676(net1979,net1981_c1,net1980_c1);
SPLITT SplitCLK_6_677(net1962,net1978_c1,net1979_c1);
SPLITT SplitCLK_6_678(net1972,net1976_c1,net1977_c1);
SPLITT SplitCLK_4_679(net1973,net1974_c1,net1975_c1);
SPLITT SplitCLK_4_680(net1964,net1972_c1,net1973_c1);
SPLITT SplitCLK_0_681(net1966,net1970_c1,net1971_c1);
SPLITT SplitCLK_2_682(net1967,net1968_c1,net1969_c1);
SPLITT SplitCLK_2_683(net1965,net1966_c1,net1967_c1);
SPLITT SplitCLK_4_684(net1963,net1965_c1,net1964_c1);
SPLITT SplitCLK_2_685(net1961,net1963_c1,net1962_c1);
SPLITT SplitCLK_6_686(net1894,net1960_c1,net1961_c1);
SPLITT SplitCLK_4_687(net1957,net1959_c1,net1958_c1);
SPLITT SplitCLK_0_688(net1952,net1956_c1,net1957_c1);
SPLITT SplitCLK_2_689(net1953,net1955_c1,net1954_c1);
SPLITT SplitCLK_4_690(net1944,net1953_c1,net1952_c1);
SPLITT SplitCLK_6_691(net1946,net1950_c1,net1951_c1);
SPLITT SplitCLK_2_692(net1947,net1948_c1,net1949_c1);
SPLITT SplitCLK_6_693(net1945,net1946_c1,net1947_c1);
SPLITT SplitCLK_4_694(net1928,net1945_c1,net1944_c1);
SPLITT SplitCLK_0_695(net1938,net1943_c1,net1942_c1);
SPLITT SplitCLK_4_696(net1939,net1941_c1,net1940_c1);
SPLITT SplitCLK_4_697(net1930,net1939_c1,net1938_c1);
SPLITT SplitCLK_6_698(net1932,net1937_c1,net1936_c1);
SPLITT SplitCLK_4_699(net1933,net1934_c1,net1935_c1);
SPLITT SplitCLK_2_700(net1931,net1933_c1,net1932_c1);
SPLITT SplitCLK_4_701(net1929,net1931_c1,net1930_c1);
SPLITT SplitCLK_0_702(net1896,net1928_c1,net1929_c1);
SPLITT SplitCLK_4_703(net1922,net1926_c1,net1927_c1);
SPLITT SplitCLK_4_704(net1923,net1925_c1,net1924_c1);
SPLITT SplitCLK_0_705(net1914,net1922_c1,net1923_c1);
SPLITT SplitCLK_6_706(net1916,net1921_c1,net1920_c1);
SPLITT SplitCLK_4_707(net1917,net1918_c1,net1919_c1);
SPLITT SplitCLK_2_708(net1915,net1917_c1,net1916_c1);
SPLITT SplitCLK_6_709(net1898,net1914_c1,net1915_c1);
SPLITT SplitCLK_4_710(net1908,net1912_c1,net1913_c1);
SPLITT SplitCLK_4_711(net1909,net1910_c1,net1911_c1);
SPLITT SplitCLK_0_712(net1900,net1908_c1,net1909_c1);
SPLITT SplitCLK_6_713(net1902,net1907_c1,net1906_c1);
SPLITT SplitCLK_6_714(net1903,net1905_c1,net1904_c1);
SPLITT SplitCLK_4_715(net1901,net1903_c1,net1902_c1);
SPLITT SplitCLK_4_716(net1899,net1901_c1,net1900_c1);
SPLITT SplitCLK_4_717(net1897,net1899_c1,net1898_c1);
SPLITT SplitCLK_4_718(net1895,net1897_c1,net1896_c1);
SPLITT SplitCLK_0_719(net1764,net1894_c1,net1895_c1);
SPLITT SplitCLK_4_720(net1891,net1893_c1,net1892_c1);
SPLITT SplitCLK_4_721(net1886,net1890_c1,net1891_c1);
SPLITT SplitCLK_4_722(net1887,net1889_c1,net1888_c1);
SPLITT SplitCLK_4_723(net1878,net1887_c1,net1886_c1);
SPLITT SplitCLK_6_724(net1880,net1885_c1,net1884_c1);
SPLITT SplitCLK_4_725(net1881,net1883_c1,net1882_c1);
SPLITT SplitCLK_6_726(net1879,net1881_c1,net1880_c1);
SPLITT SplitCLK_6_727(net1862,net1878_c1,net1879_c1);
SPLITT SplitCLK_0_728(net1872,net1877_c1,net1876_c1);
SPLITT SplitCLK_4_729(net1873,net1874_c1,net1875_c1);
SPLITT SplitCLK_4_730(net1864,net1873_c1,net1872_c1);
SPLITT SplitCLK_2_731(net1866,net1871_c1,net1870_c1);
SPLITT SplitCLK_4_732(net1867,net1869_c1,net1868_c1);
SPLITT SplitCLK_2_733(net1865,net1867_c1,net1866_c1);
SPLITT SplitCLK_4_734(net1863,net1865_c1,net1864_c1);
SPLITT SplitCLK_0_735(net1830,net1862_c1,net1863_c1);
SPLITT SplitCLK_6_736(net1856,net1860_c1,net1861_c1);
SPLITT SplitCLK_0_737(net1857,net1859_c1,net1858_c1);
SPLITT SplitCLK_4_738(net1848,net1856_c1,net1857_c1);
SPLITT SplitCLK_6_739(net1850,net1854_c1,net1855_c1);
SPLITT SplitCLK_4_740(net1851,net1852_c1,net1853_c1);
SPLITT SplitCLK_6_741(net1849,net1851_c1,net1850_c1);
SPLITT SplitCLK_6_742(net1832,net1848_c1,net1849_c1);
SPLITT SplitCLK_4_743(net1842,net1847_c1,net1846_c1);
SPLITT SplitCLK_4_744(net1843,net1844_c1,net1845_c1);
SPLITT SplitCLK_0_745(net1834,net1842_c1,net1843_c1);
SPLITT SplitCLK_6_746(net1836,net1841_c1,net1840_c1);
SPLITT SplitCLK_4_747(net1837,net1839_c1,net1838_c1);
SPLITT SplitCLK_2_748(net1835,net1836_c1,net1837_c1);
SPLITT SplitCLK_4_749(net1833,net1835_c1,net1834_c1);
SPLITT SplitCLK_2_750(net1831,net1833_c1,net1832_c1);
SPLITT SplitCLK_6_751(net1766,net1830_c1,net1831_c1);
SPLITT SplitCLK_4_752(net1824,net1828_c1,net1829_c1);
SPLITT SplitCLK_4_753(net1825,net1826_c1,net1827_c1);
SPLITT SplitCLK_0_754(net1816,net1824_c1,net1825_c1);
SPLITT SplitCLK_6_755(net1818,net1822_c1,net1823_c1);
SPLITT SplitCLK_6_756(net1819,net1821_c1,net1820_c1);
SPLITT SplitCLK_4_757(net1817,net1819_c1,net1818_c1);
SPLITT SplitCLK_6_758(net1800,net1816_c1,net1817_c1);
SPLITT SplitCLK_4_759(net1810,net1814_c1,net1815_c1);
SPLITT SplitCLK_4_760(net1811,net1812_c1,net1813_c1);
SPLITT SplitCLK_0_761(net1802,net1810_c1,net1811_c1);
SPLITT SplitCLK_6_762(net1804,net1809_c1,net1808_c1);
SPLITT SplitCLK_6_763(net1805,net1807_c1,net1806_c1);
SPLITT SplitCLK_4_764(net1803,net1805_c1,net1804_c1);
SPLITT SplitCLK_4_765(net1801,net1803_c1,net1802_c1);
SPLITT SplitCLK_0_766(net1768,net1800_c1,net1801_c1);
SPLITT SplitCLK_4_767(net1794,net1798_c1,net1799_c1);
SPLITT SplitCLK_4_768(net1795,net1796_c1,net1797_c1);
SPLITT SplitCLK_6_769(net1786,net1794_c1,net1795_c1);
SPLITT SplitCLK_6_770(net1788,net1792_c1,net1793_c1);
SPLITT SplitCLK_6_771(net1789,net1791_c1,net1790_c1);
SPLITT SplitCLK_6_772(net1787,net1788_c1,net1789_c1);
SPLITT SplitCLK_4_773(net1770,net1787_c1,net1786_c1);
SPLITT SplitCLK_4_774(net1780,net1784_c1,net1785_c1);
SPLITT SplitCLK_4_775(net1781,net1782_c1,net1783_c1);
SPLITT SplitCLK_0_776(net1772,net1780_c1,net1781_c1);
SPLITT SplitCLK_6_777(net1774,net1779_c1,net1778_c1);
SPLITT SplitCLK_4_778(net1775,net1776_c1,net1777_c1);
SPLITT SplitCLK_2_779(net1773,net1775_c1,net1774_c1);
SPLITT SplitCLK_4_780(net1771,net1773_c1,net1772_c1);
SPLITT SplitCLK_6_781(net1769,net1770_c1,net1771_c1);
SPLITT SplitCLK_4_782(net1767,net1769_c1,net1768_c1);
SPLITT SplitCLK_4_783(net1765,net1766_c1,net1767_c1);
SPLITT SplitCLK_4_784(net1763,net1765_c1,net1764_c1);
SPLITT SplitCLK_0_785(net738,net1762_c1,net1763_c1);
SPLITT SplitCLK_4_786(net1759,net1761_c1,net1760_c1);
SPLITT SplitCLK_2_787(net1754,net1758_c1,net1759_c1);
SPLITT SplitCLK_2_788(net1755,net1757_c1,net1756_c1);
SPLITT SplitCLK_4_789(net1746,net1755_c1,net1754_c1);
SPLITT SplitCLK_6_790(net1748,net1752_c1,net1753_c1);
SPLITT SplitCLK_6_791(net1749,net1750_c1,net1751_c1);
SPLITT SplitCLK_6_792(net1747,net1748_c1,net1749_c1);
SPLITT SplitCLK_6_793(net1730,net1746_c1,net1747_c1);
SPLITT SplitCLK_4_794(net1740,net1744_c1,net1745_c1);
SPLITT SplitCLK_4_795(net1741,net1743_c1,net1742_c1);
SPLITT SplitCLK_0_796(net1732,net1740_c1,net1741_c1);
SPLITT SplitCLK_6_797(net1734,net1738_c1,net1739_c1);
SPLITT SplitCLK_4_798(net1735,net1736_c1,net1737_c1);
SPLITT SplitCLK_2_799(net1733,net1735_c1,net1734_c1);
SPLITT SplitCLK_4_800(net1731,net1733_c1,net1732_c1);
SPLITT SplitCLK_0_801(net1698,net1730_c1,net1731_c1);
SPLITT SplitCLK_6_802(net1724,net1728_c1,net1729_c1);
SPLITT SplitCLK_0_803(net1725,net1727_c1,net1726_c1);
SPLITT SplitCLK_0_804(net1716,net1724_c1,net1725_c1);
SPLITT SplitCLK_6_805(net1718,net1722_c1,net1723_c1);
SPLITT SplitCLK_6_806(net1719,net1720_c1,net1721_c1);
SPLITT SplitCLK_6_807(net1717,net1718_c1,net1719_c1);
SPLITT SplitCLK_6_808(net1700,net1716_c1,net1717_c1);
SPLITT SplitCLK_6_809(net1710,net1714_c1,net1715_c1);
SPLITT SplitCLK_4_810(net1711,net1712_c1,net1713_c1);
SPLITT SplitCLK_4_811(net1702,net1710_c1,net1711_c1);
SPLITT SplitCLK_6_812(net1704,net1709_c1,net1708_c1);
SPLITT SplitCLK_4_813(net1705,net1707_c1,net1706_c1);
SPLITT SplitCLK_2_814(net1703,net1705_c1,net1704_c1);
SPLITT SplitCLK_4_815(net1701,net1703_c1,net1702_c1);
SPLITT SplitCLK_2_816(net1699,net1701_c1,net1700_c1);
SPLITT SplitCLK_6_817(net1632,net1698_c1,net1699_c1);
SPLITT SplitCLK_4_818(net1695,net1696_c1,net1697_c1);
SPLITT SplitCLK_2_819(net1690,net1694_c1,net1695_c1);
SPLITT SplitCLK_4_820(net1691,net1693_c1,net1692_c1);
SPLITT SplitCLK_0_821(net1682,net1690_c1,net1691_c1);
SPLITT SplitCLK_4_822(net1684,net1689_c1,net1688_c1);
SPLITT SplitCLK_4_823(net1685,net1687_c1,net1686_c1);
SPLITT SplitCLK_6_824(net1683,net1684_c1,net1685_c1);
SPLITT SplitCLK_4_825(net1666,net1683_c1,net1682_c1);
SPLITT SplitCLK_4_826(net1676,net1680_c1,net1681_c1);
SPLITT SplitCLK_4_827(net1677,net1678_c1,net1679_c1);
SPLITT SplitCLK_0_828(net1668,net1676_c1,net1677_c1);
SPLITT SplitCLK_6_829(net1670,net1675_c1,net1674_c1);
SPLITT SplitCLK_4_830(net1671,net1672_c1,net1673_c1);
SPLITT SplitCLK_2_831(net1669,net1671_c1,net1670_c1);
SPLITT SplitCLK_4_832(net1667,net1669_c1,net1668_c1);
SPLITT SplitCLK_0_833(net1634,net1666_c1,net1667_c1);
SPLITT SplitCLK_6_834(net1660,net1664_c1,net1665_c1);
SPLITT SplitCLK_4_835(net1661,net1662_c1,net1663_c1);
SPLITT SplitCLK_0_836(net1652,net1660_c1,net1661_c1);
SPLITT SplitCLK_2_837(net1654,net1658_c1,net1659_c1);
SPLITT SplitCLK_4_838(net1655,net1657_c1,net1656_c1);
SPLITT SplitCLK_6_839(net1653,net1655_c1,net1654_c1);
SPLITT SplitCLK_6_840(net1636,net1652_c1,net1653_c1);
SPLITT SplitCLK_6_841(net1646,net1651_c1,net1650_c1);
SPLITT SplitCLK_4_842(net1647,net1648_c1,net1649_c1);
SPLITT SplitCLK_0_843(net1638,net1646_c1,net1647_c1);
SPLITT SplitCLK_6_844(net1640,net1644_c1,net1645_c1);
SPLITT SplitCLK_4_845(net1641,net1642_c1,net1643_c1);
SPLITT SplitCLK_6_846(net1639,net1640_c1,net1641_c1);
SPLITT SplitCLK_4_847(net1637,net1639_c1,net1638_c1);
SPLITT SplitCLK_4_848(net1635,net1636_c1,net1637_c1);
SPLITT SplitCLK_4_849(net1633,net1635_c1,net1634_c1);
SPLITT SplitCLK_6_850(net1502,net1633_c1,net1632_c1);
SPLITT SplitCLK_4_851(net1629,net1631_c1,net1630_c1);
SPLITT SplitCLK_4_852(net1624,net1628_c1,net1629_c1);
SPLITT SplitCLK_4_853(net1625,net1627_c1,net1626_c1);
SPLITT SplitCLK_6_854(net1616,net1624_c1,net1625_c1);
SPLITT SplitCLK_6_855(net1618,net1622_c1,net1623_c1);
SPLITT SplitCLK_0_856(net1619,net1621_c1,net1620_c1);
SPLITT SplitCLK_2_857(net1617,net1619_c1,net1618_c1);
SPLITT SplitCLK_6_858(net1600,net1616_c1,net1617_c1);
SPLITT SplitCLK_6_859(net1610,net1614_c1,net1615_c1);
SPLITT SplitCLK_4_860(net1611,net1613_c1,net1612_c1);
SPLITT SplitCLK_4_861(net1602,net1611_c1,net1610_c1);
SPLITT SplitCLK_4_862(net1604,net1609_c1,net1608_c1);
SPLITT SplitCLK_6_863(net1605,net1606_c1,net1607_c1);
SPLITT SplitCLK_6_864(net1603,net1604_c1,net1605_c1);
SPLITT SplitCLK_4_865(net1601,net1603_c1,net1602_c1);
SPLITT SplitCLK_0_866(net1568,net1600_c1,net1601_c1);
SPLITT SplitCLK_6_867(net1594,net1598_c1,net1599_c1);
SPLITT SplitCLK_0_868(net1595,net1597_c1,net1596_c1);
SPLITT SplitCLK_0_869(net1586,net1594_c1,net1595_c1);
SPLITT SplitCLK_6_870(net1588,net1592_c1,net1593_c1);
SPLITT SplitCLK_4_871(net1589,net1591_c1,net1590_c1);
SPLITT SplitCLK_6_872(net1587,net1589_c1,net1588_c1);
SPLITT SplitCLK_6_873(net1570,net1586_c1,net1587_c1);
SPLITT SplitCLK_6_874(net1580,net1584_c1,net1585_c1);
SPLITT SplitCLK_0_875(net1581,net1582_c1,net1583_c1);
SPLITT SplitCLK_4_876(net1572,net1581_c1,net1580_c1);
SPLITT SplitCLK_0_877(net1574,net1578_c1,net1579_c1);
SPLITT SplitCLK_0_878(net1575,net1577_c1,net1576_c1);
SPLITT SplitCLK_2_879(net1573,net1575_c1,net1574_c1);
SPLITT SplitCLK_4_880(net1571,net1573_c1,net1572_c1);
SPLITT SplitCLK_2_881(net1569,net1571_c1,net1570_c1);
SPLITT SplitCLK_6_882(net1504,net1568_c1,net1569_c1);
SPLITT SplitCLK_0_883(net1562,net1567_c1,net1566_c1);
SPLITT SplitCLK_4_884(net1563,net1565_c1,net1564_c1);
SPLITT SplitCLK_4_885(net1554,net1562_c1,net1563_c1);
SPLITT SplitCLK_6_886(net1556,net1560_c1,net1561_c1);
SPLITT SplitCLK_4_887(net1557,net1559_c1,net1558_c1);
SPLITT SplitCLK_2_888(net1555,net1557_c1,net1556_c1);
SPLITT SplitCLK_6_889(net1538,net1554_c1,net1555_c1);
SPLITT SplitCLK_6_890(net1548,net1552_c1,net1553_c1);
SPLITT SplitCLK_0_891(net1549,net1550_c1,net1551_c1);
SPLITT SplitCLK_0_892(net1540,net1548_c1,net1549_c1);
SPLITT SplitCLK_2_893(net1542,net1546_c1,net1547_c1);
SPLITT SplitCLK_4_894(net1543,net1544_c1,net1545_c1);
SPLITT SplitCLK_6_895(net1541,net1543_c1,net1542_c1);
SPLITT SplitCLK_4_896(net1539,net1541_c1,net1540_c1);
SPLITT SplitCLK_0_897(net1506,net1538_c1,net1539_c1);
SPLITT SplitCLK_0_898(net1532,net1537_c1,net1536_c1);
SPLITT SplitCLK_4_899(net1533,net1535_c1,net1534_c1);
SPLITT SplitCLK_0_900(net1524,net1532_c1,net1533_c1);
SPLITT SplitCLK_6_901(net1526,net1531_c1,net1530_c1);
SPLITT SplitCLK_4_902(net1527,net1528_c1,net1529_c1);
SPLITT SplitCLK_6_903(net1525,net1527_c1,net1526_c1);
SPLITT SplitCLK_6_904(net1508,net1524_c1,net1525_c1);
SPLITT SplitCLK_0_905(net1518,net1523_c1,net1522_c1);
SPLITT SplitCLK_4_906(net1519,net1521_c1,net1520_c1);
SPLITT SplitCLK_4_907(net1510,net1518_c1,net1519_c1);
SPLITT SplitCLK_6_908(net1512,net1516_c1,net1517_c1);
SPLITT SplitCLK_4_909(net1513,net1515_c1,net1514_c1);
SPLITT SplitCLK_2_910(net1511,net1513_c1,net1512_c1);
SPLITT SplitCLK_4_911(net1509,net1511_c1,net1510_c1);
SPLITT SplitCLK_2_912(net1507,net1509_c1,net1508_c1);
SPLITT SplitCLK_4_913(net1505,net1507_c1,net1506_c1);
SPLITT SplitCLK_2_914(net1503,net1505_c1,net1504_c1);
SPLITT SplitCLK_6_915(net1240,net1502_c1,net1503_c1);
SPLITT SplitCLK_4_916(net1499,net1501_c1,net1500_c1);
SPLITT SplitCLK_4_917(net1494,net1498_c1,net1499_c1);
SPLITT SplitCLK_4_918(net1495,net1497_c1,net1496_c1);
SPLITT SplitCLK_6_919(net1486,net1494_c1,net1495_c1);
SPLITT SplitCLK_6_920(net1488,net1493_c1,net1492_c1);
SPLITT SplitCLK_4_921(net1489,net1491_c1,net1490_c1);
SPLITT SplitCLK_2_922(net1487,net1489_c1,net1488_c1);
SPLITT SplitCLK_6_923(net1470,net1486_c1,net1487_c1);
SPLITT SplitCLK_6_924(net1480,net1485_c1,net1484_c1);
SPLITT SplitCLK_0_925(net1481,net1482_c1,net1483_c1);
SPLITT SplitCLK_0_926(net1472,net1480_c1,net1481_c1);
SPLITT SplitCLK_0_927(net1474,net1478_c1,net1479_c1);
SPLITT SplitCLK_6_928(net1475,net1476_c1,net1477_c1);
SPLITT SplitCLK_6_929(net1473,net1474_c1,net1475_c1);
SPLITT SplitCLK_4_930(net1471,net1473_c1,net1472_c1);
SPLITT SplitCLK_0_931(net1438,net1470_c1,net1471_c1);
SPLITT SplitCLK_0_932(net1464,net1468_c1,net1469_c1);
SPLITT SplitCLK_2_933(net1465,net1467_c1,net1466_c1);
SPLITT SplitCLK_4_934(net1456,net1465_c1,net1464_c1);
SPLITT SplitCLK_6_935(net1458,net1462_c1,net1463_c1);
SPLITT SplitCLK_4_936(net1459,net1461_c1,net1460_c1);
SPLITT SplitCLK_2_937(net1457,net1459_c1,net1458_c1);
SPLITT SplitCLK_6_938(net1440,net1456_c1,net1457_c1);
SPLITT SplitCLK_6_939(net1450,net1454_c1,net1455_c1);
SPLITT SplitCLK_4_940(net1451,net1453_c1,net1452_c1);
SPLITT SplitCLK_4_941(net1442,net1450_c1,net1451_c1);
SPLITT SplitCLK_0_942(net1444,net1449_c1,net1448_c1);
SPLITT SplitCLK_6_943(net1445,net1447_c1,net1446_c1);
SPLITT SplitCLK_6_944(net1443,net1444_c1,net1445_c1);
SPLITT SplitCLK_4_945(net1441,net1443_c1,net1442_c1);
SPLITT SplitCLK_2_946(net1439,net1441_c1,net1440_c1);
SPLITT SplitCLK_6_947(net1372,net1438_c1,net1439_c1);
SPLITT SplitCLK_4_948(net1435,net1436_c1,net1437_c1);
SPLITT SplitCLK_0_949(net1430,net1434_c1,net1435_c1);
SPLITT SplitCLK_0_950(net1431,net1432_c1,net1433_c1);
SPLITT SplitCLK_4_951(net1422,net1430_c1,net1431_c1);
SPLITT SplitCLK_0_952(net1424,net1429_c1,net1428_c1);
SPLITT SplitCLK_4_953(net1425,net1427_c1,net1426_c1);
SPLITT SplitCLK_2_954(net1423,net1425_c1,net1424_c1);
SPLITT SplitCLK_6_955(net1406,net1422_c1,net1423_c1);
SPLITT SplitCLK_6_956(net1416,net1420_c1,net1421_c1);
SPLITT SplitCLK_4_957(net1417,net1418_c1,net1419_c1);
SPLITT SplitCLK_0_958(net1408,net1416_c1,net1417_c1);
SPLITT SplitCLK_6_959(net1410,net1414_c1,net1415_c1);
SPLITT SplitCLK_6_960(net1411,net1412_c1,net1413_c1);
SPLITT SplitCLK_6_961(net1409,net1410_c1,net1411_c1);
SPLITT SplitCLK_4_962(net1407,net1409_c1,net1408_c1);
SPLITT SplitCLK_0_963(net1374,net1406_c1,net1407_c1);
SPLITT SplitCLK_4_964(net1400,net1405_c1,net1404_c1);
SPLITT SplitCLK_4_965(net1401,net1403_c1,net1402_c1);
SPLITT SplitCLK_6_966(net1392,net1400_c1,net1401_c1);
SPLITT SplitCLK_6_967(net1394,net1399_c1,net1398_c1);
SPLITT SplitCLK_6_968(net1395,net1396_c1,net1397_c1);
SPLITT SplitCLK_6_969(net1393,net1394_c1,net1395_c1);
SPLITT SplitCLK_6_970(net1376,net1392_c1,net1393_c1);
SPLITT SplitCLK_4_971(net1386,net1390_c1,net1391_c1);
SPLITT SplitCLK_4_972(net1387,net1388_c1,net1389_c1);
SPLITT SplitCLK_4_973(net1378,net1387_c1,net1386_c1);
SPLITT SplitCLK_6_974(net1380,net1384_c1,net1385_c1);
SPLITT SplitCLK_4_975(net1381,net1383_c1,net1382_c1);
SPLITT SplitCLK_2_976(net1379,net1381_c1,net1380_c1);
SPLITT SplitCLK_4_977(net1377,net1379_c1,net1378_c1);
SPLITT SplitCLK_2_978(net1375,net1377_c1,net1376_c1);
SPLITT SplitCLK_4_979(net1373,net1375_c1,net1374_c1);
SPLITT SplitCLK_0_980(net1242,net1372_c1,net1373_c1);
SPLITT SplitCLK_4_981(net1369,net1370_c1,net1371_c1);
SPLITT SplitCLK_4_982(net1364,net1368_c1,net1369_c1);
SPLITT SplitCLK_4_983(net1365,net1366_c1,net1367_c1);
SPLITT SplitCLK_0_984(net1356,net1364_c1,net1365_c1);
SPLITT SplitCLK_6_985(net1358,net1363_c1,net1362_c1);
SPLITT SplitCLK_0_986(net1359,net1360_c1,net1361_c1);
SPLITT SplitCLK_6_987(net1357,net1359_c1,net1358_c1);
SPLITT SplitCLK_6_988(net1340,net1356_c1,net1357_c1);
SPLITT SplitCLK_4_989(net1350,net1354_c1,net1355_c1);
SPLITT SplitCLK_4_990(net1351,net1352_c1,net1353_c1);
SPLITT SplitCLK_6_991(net1342,net1350_c1,net1351_c1);
SPLITT SplitCLK_0_992(net1344,net1348_c1,net1349_c1);
SPLITT SplitCLK_6_993(net1345,net1347_c1,net1346_c1);
SPLITT SplitCLK_6_994(net1343,net1344_c1,net1345_c1);
SPLITT SplitCLK_4_995(net1341,net1343_c1,net1342_c1);
SPLITT SplitCLK_0_996(net1308,net1340_c1,net1341_c1);
SPLITT SplitCLK_0_997(net1334,net1339_c1,net1338_c1);
SPLITT SplitCLK_0_998(net1335,net1337_c1,net1336_c1);
SPLITT SplitCLK_2_999(net1326,net1335_c1,net1334_c1);
SPLITT SplitCLK_6_1000(net1328,net1333_c1,net1332_c1);
SPLITT SplitCLK_4_1001(net1329,net1331_c1,net1330_c1);
SPLITT SplitCLK_6_1002(net1327,net1328_c1,net1329_c1);
SPLITT SplitCLK_6_1003(net1310,net1326_c1,net1327_c1);
SPLITT SplitCLK_0_1004(net1320,net1324_c1,net1325_c1);
SPLITT SplitCLK_4_1005(net1321,net1323_c1,net1322_c1);
SPLITT SplitCLK_4_1006(net1312,net1321_c1,net1320_c1);
SPLITT SplitCLK_6_1007(net1314,net1318_c1,net1319_c1);
SPLITT SplitCLK_4_1008(net1315,net1316_c1,net1317_c1);
SPLITT SplitCLK_6_1009(net1313,net1314_c1,net1315_c1);
SPLITT SplitCLK_4_1010(net1311,net1313_c1,net1312_c1);
SPLITT SplitCLK_4_1011(net1309,net1310_c1,net1311_c1);
SPLITT SplitCLK_6_1012(net1244,net1308_c1,net1309_c1);
SPLITT SplitCLK_0_1013(net1302,net1307_c1,net1306_c1);
SPLITT SplitCLK_2_1014(net1303,net1305_c1,net1304_c1);
SPLITT SplitCLK_4_1015(net1294,net1303_c1,net1302_c1);
SPLITT SplitCLK_6_1016(net1296,net1300_c1,net1301_c1);
SPLITT SplitCLK_4_1017(net1297,net1298_c1,net1299_c1);
SPLITT SplitCLK_2_1018(net1295,net1297_c1,net1296_c1);
SPLITT SplitCLK_6_1019(net1278,net1294_c1,net1295_c1);
SPLITT SplitCLK_6_1020(net1288,net1292_c1,net1293_c1);
SPLITT SplitCLK_4_1021(net1289,net1291_c1,net1290_c1);
SPLITT SplitCLK_0_1022(net1280,net1288_c1,net1289_c1);
SPLITT SplitCLK_0_1023(net1282,net1287_c1,net1286_c1);
SPLITT SplitCLK_6_1024(net1283,net1284_c1,net1285_c1);
SPLITT SplitCLK_2_1025(net1281,net1282_c1,net1283_c1);
SPLITT SplitCLK_4_1026(net1279,net1281_c1,net1280_c1);
SPLITT SplitCLK_0_1027(net1246,net1278_c1,net1279_c1);
SPLITT SplitCLK_6_1028(net1272,net1277_c1,net1276_c1);
SPLITT SplitCLK_4_1029(net1273,net1275_c1,net1274_c1);
SPLITT SplitCLK_0_1030(net1264,net1272_c1,net1273_c1);
SPLITT SplitCLK_6_1031(net1266,net1271_c1,net1270_c1);
SPLITT SplitCLK_4_1032(net1267,net1269_c1,net1268_c1);
SPLITT SplitCLK_6_1033(net1265,net1267_c1,net1266_c1);
SPLITT SplitCLK_6_1034(net1248,net1264_c1,net1265_c1);
SPLITT SplitCLK_4_1035(net1258,net1263_c1,net1262_c1);
SPLITT SplitCLK_4_1036(net1259,net1260_c1,net1261_c1);
SPLITT SplitCLK_4_1037(net1250,net1259_c1,net1258_c1);
SPLITT SplitCLK_6_1038(net1252,net1256_c1,net1257_c1);
SPLITT SplitCLK_4_1039(net1253,net1254_c1,net1255_c1);
SPLITT SplitCLK_2_1040(net1251,net1253_c1,net1252_c1);
SPLITT SplitCLK_4_1041(net1249,net1251_c1,net1250_c1);
SPLITT SplitCLK_2_1042(net1247,net1249_c1,net1248_c1);
SPLITT SplitCLK_4_1043(net1245,net1247_c1,net1246_c1);
SPLITT SplitCLK_2_1044(net1243,net1245_c1,net1244_c1);
SPLITT SplitCLK_4_1045(net1241,net1243_c1,net1242_c1);
SPLITT SplitCLK_2_1046(net739,net1241_c1,net1240_c1);
wire dummy0;
SPLITT SplitCLK_4_1047(net1722,net1239_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_4_1048(net2014,net1238_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_4_1049(net1940,net1237_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_1050(net1812,net1236_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_1051(net2018,net1235_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_2_1052(net1426,net1234_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_4_1053(net1262,net1233_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_4_1054(net1336,net1232_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_4_1055(net1838,net1231_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_4_1056(net1664,net1230_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_2_1057(net1796,net1229_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_2_1058(net1530,net1228_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_4_1059(net2264,net1227_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_4_1060(net1598,net1226_c1,dummy13);
wire dummy14;
SPLITT SplitCLK_2_1061(net1723,net1225_c1,dummy14);
wire dummy15;
SPLITT SplitCLK_2_1062(net2150,net1224_c1,dummy15);
wire dummy16;
SPLITT SplitCLK_4_1063(net1558,net1223_c1,dummy16);
wire dummy17;
SPLITT SplitCLK_4_1064(net2012,net1222_c1,dummy17);
wire dummy18;
SPLITT SplitCLK_2_1065(net2202,net1221_c1,dummy18);
wire dummy19;
SPLITT SplitCLK_2_1066(net1941,net1220_c1,dummy19);
wire dummy20;
SPLITT SplitCLK_4_1067(net1813,net1219_c1,dummy20);
wire dummy21;
SPLITT SplitCLK_4_1068(net1792,net1218_c1,dummy21);
wire dummy22;
SPLITT SplitCLK_4_1069(net1428,net1217_c1,dummy22);
wire dummy23;
SPLITT SplitCLK_2_1070(net1263,net1216_c1,dummy23);
wire dummy24;
SPLITT SplitCLK_2_1071(net1354,net1215_c1,dummy24);
wire dummy25;
SPLITT SplitCLK_4_1072(net1644,net1214_c1,dummy25);
wire dummy26;
SPLITT SplitCLK_4_1073(net1797,net1213_c1,dummy26);
wire dummy27;
SPLITT SplitCLK_4_1074(net2144,net1212_c1,dummy27);
wire dummy28;
SPLITT SplitCLK_4_1075(net1536,net1211_c1,dummy28);
wire dummy29;
SPLITT SplitCLK_4_1076(net2006,net1210_c1,dummy29);
wire dummy30;
SPLITT SplitCLK_4_1077(net2203,net1209_c1,dummy30);
wire dummy31;
SPLITT SplitCLK_4_1078(net1942,net1208_c1,dummy31);
wire dummy32;
SPLITT SplitCLK_2_1079(net1904,net1207_c1,dummy32);
wire dummy33;
SPLITT SplitCLK_2_1080(net1348,net1206_c1,dummy33);
wire dummy34;
SPLITT SplitCLK_2_1081(net1432,net1205_c1,dummy34);
wire dummy35;
SPLITT SplitCLK_2_1082(net1260,net1204_c1,dummy35);
wire dummy36;
SPLITT SplitCLK_2_1083(net1388,net1203_c1,dummy36);
wire dummy37;
SPLITT SplitCLK_4_1084(net1656,net1202_c1,dummy37);
wire dummy38;
SPLITT SplitCLK_2_1085(net1820,net1201_c1,dummy38);
wire dummy39;
SPLITT SplitCLK_4_1086(net1821,net1200_c1,dummy39);
wire dummy40;
SPLITT SplitCLK_4_1087(net1414,net1199_c1,dummy40);
wire dummy41;
SPLITT SplitCLK_4_1088(net2004,net1198_c1,dummy41);
wire dummy42;
SPLITT SplitCLK_2_1089(net2196,net1197_c1,dummy42);
wire dummy43;
SPLITT SplitCLK_4_1090(net1943,net1196_c1,dummy43);
wire dummy44;
SPLITT SplitCLK_4_1091(net1349,net1195_c1,dummy44);
wire dummy45;
SPLITT SplitCLK_2_1092(net1490,net1194_c1,dummy45);
wire dummy46;
SPLITT SplitCLK_4_1093(net1256,net1193_c1,dummy46);
wire dummy47;
SPLITT SplitCLK_2_1094(net1650,net1192_c1,dummy47);
wire dummy48;
SPLITT SplitCLK_2_1095(net1706,net1191_c1,dummy48);
wire dummy49;
SPLITT SplitCLK_2_1096(net2250,net1190_c1,dummy49);
wire dummy50;
SPLITT SplitCLK_2_1097(net1366,net1189_c1,dummy50);
wire dummy51;
SPLITT SplitCLK_4_1098(net2128,net1188_c1,dummy51);
wire dummy52;
SPLITT SplitCLK_4_1099(net2265,net1187_c1,dummy52);
wire dummy53;
SPLITT SplitCLK_4_1100(net1714,net1186_c1,dummy53);
wire dummy54;
SPLITT SplitCLK_2_1101(net1688,net1185_c1,dummy54);
wire dummy55;
SPLITT SplitCLK_2_1102(net1537,net1184_c1,dummy55);
wire dummy56;
SPLITT SplitCLK_2_1103(net1954,net1183_c1,dummy56);
wire dummy57;
SPLITT SplitCLK_2_1104(net1852,net1182_c1,dummy57);
wire dummy58;
SPLITT SplitCLK_4_1105(net1318,net1181_c1,dummy58);
wire dummy59;
SPLITT SplitCLK_4_1106(net2044,net1180_c1,dummy59);
wire dummy60;
SPLITT SplitCLK_4_1107(net1982,net1179_c1,dummy60);
wire dummy61;
SPLITT SplitCLK_4_1108(net1346,net1178_c1,dummy61);
wire dummy62;
SPLITT SplitCLK_4_1109(net1686,net1177_c1,dummy62);
wire dummy63;
SPLITT SplitCLK_4_1110(net1988,net1176_c1,dummy63);
wire dummy64;
SPLITT SplitCLK_4_1111(net1306,net1175_c1,dummy64);
wire dummy65;
SPLITT SplitCLK_4_1112(net1404,net1174_c1,dummy65);
wire dummy66;
SPLITT SplitCLK_2_1113(net1492,net1173_c1,dummy66);
wire dummy67;
SPLITT SplitCLK_2_1114(net1926,net1172_c1,dummy67);
wire dummy68;
SPLITT SplitCLK_2_1115(net1276,net1171_c1,dummy68);
wire dummy69;
SPLITT SplitCLK_2_1116(net1478,net1170_c1,dummy69);
wire dummy70;
SPLITT SplitCLK_4_1117(net1882,net1169_c1,dummy70);
wire dummy71;
SPLITT SplitCLK_2_1118(net2244,net1168_c1,dummy71);
wire dummy72;
SPLITT SplitCLK_2_1119(net1826,net1167_c1,dummy72);
wire dummy73;
SPLITT SplitCLK_4_1120(net1420,net1166_c1,dummy73);
wire dummy74;
SPLITT SplitCLK_2_1121(net2005,net1165_c1,dummy74);
wire dummy75;
SPLITT SplitCLK_2_1122(net2200,net1164_c1,dummy75);
wire dummy76;
SPLITT SplitCLK_4_1123(net1955,net1163_c1,dummy76);
wire dummy77;
SPLITT SplitCLK_4_1124(net1347,net1162_c1,dummy77);
wire dummy78;
SPLITT SplitCLK_4_1125(net1479,net1161_c1,dummy78);
wire dummy79;
SPLITT SplitCLK_2_1126(net1257,net1160_c1,dummy79);
wire dummy80;
SPLITT SplitCLK_2_1127(net1657,net1159_c1,dummy80);
wire dummy81;
SPLITT SplitCLK_4_1128(net1827,net1158_c1,dummy81);
wire dummy82;
SPLITT SplitCLK_2_1129(net1778,net1157_c1,dummy82);
wire dummy83;
SPLITT SplitCLK_2_1130(net1956,net1156_c1,dummy83);
wire dummy84;
SPLITT SplitCLK_4_1131(net2201,net1155_c1,dummy84);
wire dummy85;
SPLITT SplitCLK_4_1132(net1322,net1154_c1,dummy85);
wire dummy86;
SPLITT SplitCLK_2_1133(net1482,net1153_c1,dummy86);
wire dummy87;
SPLITT SplitCLK_2_1134(net1254,net1152_c1,dummy87);
wire dummy88;
SPLITT SplitCLK_2_1135(net1758,net1151_c1,dummy88);
wire dummy89;
SPLITT SplitCLK_2_1136(net2145,net1150_c1,dummy89);
wire dummy90;
SPLITT SplitCLK_2_1137(net1918,net1149_c1,dummy90);
wire dummy91;
SPLITT SplitCLK_4_1138(net1779,net1148_c1,dummy91);
wire dummy92;
SPLITT SplitCLK_4_1139(net1658,net1147_c1,dummy92);
wire dummy93;
SPLITT SplitCLK_2_1140(net1307,net1146_c1,dummy93);
wire dummy94;
SPLITT SplitCLK_2_1141(net1839,net1145_c1,dummy94);
wire dummy95;
SPLITT SplitCLK_2_1142(net1920,net1144_c1,dummy95);
wire dummy96;
SPLITT SplitCLK_2_1143(net1784,net1143_c1,dummy96);
wire dummy97;
SPLITT SplitCLK_4_1144(net1564,net1142_c1,dummy97);
wire dummy98;
SPLITT SplitCLK_4_1145(net1352,net1141_c1,dummy98);
wire dummy99;
SPLITT SplitCLK_4_1146(net1921,net1140_c1,dummy99);
wire dummy100;
SPLITT SplitCLK_4_1147(net1785,net1139_c1,dummy100);
wire dummy101;
SPLITT SplitCLK_2_1148(net1565,net1138_c1,dummy101);
wire dummy102;
SPLITT SplitCLK_2_1149(net1398,net1137_c1,dummy102);
wire dummy103;
SPLITT SplitCLK_2_1150(net1793,net1136_c1,dummy103);
wire dummy104;
SPLITT SplitCLK_2_1151(net1715,net1135_c1,dummy104);
wire dummy105;
SPLITT SplitCLK_2_1152(net1712,net1134_c1,dummy105);
wire dummy106;
SPLITT SplitCLK_4_1153(net2134,net1133_c1,dummy106);
wire dummy107;
SPLITT SplitCLK_2_1154(net2098,net1132_c1,dummy107);
wire dummy108;
SPLITT SplitCLK_4_1155(net1614,net1131_c1,dummy108);
wire dummy109;
SPLITT SplitCLK_2_1156(net1608,net1130_c1,dummy109);
wire dummy110;
SPLITT SplitCLK_2_1157(net1689,net1129_c1,dummy110);
wire dummy111;
SPLITT SplitCLK_2_1158(net1708,net1128_c1,dummy111);
wire dummy112;
SPLITT SplitCLK_4_1159(net2242,net1127_c1,dummy112);
wire dummy113;
SPLITT SplitCLK_4_1160(net1626,net1126_c1,dummy113);
wire dummy114;
SPLITT SplitCLK_2_1161(net1687,net1125_c1,dummy114);
wire dummy115;
SPLITT SplitCLK_2_1162(net1756,net1124_c1,dummy115);
wire dummy116;
SPLITT SplitCLK_4_1163(net2050,net1123_c1,dummy116);
wire dummy117;
SPLITT SplitCLK_2_1164(net2129,net1122_c1,dummy117);
wire dummy118;
SPLITT SplitCLK_2_1165(net2130,net1121_c1,dummy118);
wire dummy119;
SPLITT SplitCLK_4_1166(net2148,net1120_c1,dummy119);
wire dummy120;
SPLITT SplitCLK_2_1167(net2234,net1119_c1,dummy120);
wire dummy121;
SPLITT SplitCLK_4_1168(net1860,net1118_c1,dummy121);
wire dummy122;
SPLITT SplitCLK_4_1169(net2104,net1117_c1,dummy122);
wire dummy123;
SPLITT SplitCLK_2_1170(net2278,net1116_c1,dummy123);
wire dummy124;
SPLITT SplitCLK_4_1171(net2088,net1115_c1,dummy124);
wire dummy125;
SPLITT SplitCLK_2_1172(net2080,net1114_c1,dummy125);
wire dummy126;
SPLITT SplitCLK_2_1173(net1672,net1113_c1,dummy126);
wire dummy127;
SPLITT SplitCLK_4_1174(net2056,net1112_c1,dummy127);
wire dummy128;
SPLITT SplitCLK_4_1175(net1692,net1111_c1,dummy128);
wire dummy129;
SPLITT SplitCLK_4_1176(net1858,net1110_c1,dummy129);
wire dummy130;
SPLITT SplitCLK_2_1177(net1990,net1109_c1,dummy130);
wire dummy131;
SPLITT SplitCLK_4_1178(net1476,net1108_c1,dummy131);
wire dummy132;
SPLITT SplitCLK_2_1179(net1477,net1107_c1,dummy132);
wire dummy133;
SPLITT SplitCLK_2_1180(net1736,net1106_c1,dummy133);
wire dummy134;
SPLITT SplitCLK_4_1181(net2266,net1105_c1,dummy134);
wire dummy135;
SPLITT SplitCLK_4_1182(net1454,net1104_c1,dummy135);
wire dummy136;
SPLITT SplitCLK_2_1183(net1808,net1103_c1,dummy136);
wire dummy137;
SPLITT SplitCLK_4_1184(net2058,net1102_c1,dummy137);
wire dummy138;
SPLITT SplitCLK_2_1185(net1390,net1101_c1,dummy138);
wire dummy139;
SPLITT SplitCLK_4_1186(net1809,net1100_c1,dummy139);
wire dummy140;
SPLITT SplitCLK_4_1187(net1546,net1099_c1,dummy140);
wire dummy141;
SPLITT SplitCLK_2_1188(net2136,net1098_c1,dummy141);
wire dummy142;
SPLITT SplitCLK_4_1189(net1391,net1097_c1,dummy142);
wire dummy143;
SPLITT SplitCLK_2_1190(net2000,net1096_c1,dummy143);
wire dummy144;
SPLITT SplitCLK_4_1191(net1300,net1095_c1,dummy144);
wire dummy145;
SPLITT SplitCLK_4_1192(net1738,net1094_c1,dummy145);
wire dummy146;
SPLITT SplitCLK_2_1193(net1693,net1093_c1,dummy146);
wire dummy147;
SPLITT SplitCLK_2_1194(net1694,net1092_c1,dummy147);
wire dummy148;
SPLITT SplitCLK_4_1195(net1726,net1091_c1,dummy148);
wire dummy149;
SPLITT SplitCLK_2_1196(net1739,net1090_c1,dummy149);
wire dummy150;
SPLITT SplitCLK_2_1197(net1744,net1089_c1,dummy150);
wire dummy151;
SPLITT SplitCLK_4_1198(net1620,net1088_c1,dummy151);
wire dummy152;
SPLITT SplitCLK_2_1199(net2228,net1087_c1,dummy152);
wire dummy153;
SPLITT SplitCLK_4_1200(net1742,net1086_c1,dummy153);
wire dummy154;
SPLITT SplitCLK_2_1201(net2272,net1085_c1,dummy154);
wire dummy155;
SPLITT SplitCLK_4_1202(net2099,net1084_c1,dummy155);
wire dummy156;
SPLITT SplitCLK_2_1203(net2251,net1083_c1,dummy156);
wire dummy157;
SPLITT SplitCLK_4_1204(net1615,net1082_c1,dummy157);
wire dummy158;
SPLITT SplitCLK_2_1205(net2106,net1081_c1,dummy158);
wire dummy159;
SPLITT SplitCLK_4_1206(net1720,net1080_c1,dummy159);
wire dummy160;
SPLITT SplitCLK_4_1207(net2248,net1079_c1,dummy160);
wire dummy161;
SPLITT SplitCLK_4_1208(net1460,net1078_c1,dummy161);
wire dummy162;
SPLITT SplitCLK_4_1209(net2100,net1077_c1,dummy162);
wire dummy163;
SPLITT SplitCLK_4_1210(net1483,net1076_c1,dummy163);
wire dummy164;
SPLITT SplitCLK_2_1211(net2107,net1075_c1,dummy164);
wire dummy165;
SPLITT SplitCLK_2_1212(net2149,net1074_c1,dummy165);
wire dummy166;
SPLITT SplitCLK_4_1213(net2072,net1073_c1,dummy166);
wire dummy167;
SPLITT SplitCLK_4_1214(net1984,net1072_c1,dummy167);
wire dummy168;
SPLITT SplitCLK_2_1215(net1582,net1071_c1,dummy168);
wire dummy169;
SPLITT SplitCLK_2_1216(net1870,net1070_c1,dummy169);
wire dummy170;
SPLITT SplitCLK_4_1217(net2082,net1069_c1,dummy170);
wire dummy171;
SPLITT SplitCLK_2_1218(net1491,net1068_c1,dummy171);
wire dummy172;
SPLITT SplitCLK_2_1219(net1665,net1067_c1,dummy172);
wire dummy173;
SPLITT SplitCLK_4_1220(net1651,net1066_c1,dummy173);
wire dummy174;
SPLITT SplitCLK_2_1221(net1550,net1065_c1,dummy174);
wire dummy175;
SPLITT SplitCLK_2_1222(net2135,net1064_c1,dummy175);
wire dummy176;
SPLITT SplitCLK_4_1223(net1412,net1063_c1,dummy176);
wire dummy177;
SPLITT SplitCLK_4_1224(net1534,net1062_c1,dummy177);
wire dummy178;
SPLITT SplitCLK_4_1225(net1552,net1061_c1,dummy178);
wire dummy179;
SPLITT SplitCLK_4_1226(net1551,net1060_c1,dummy179);
wire dummy180;
SPLITT SplitCLK_2_1227(net2089,net1059_c1,dummy180);
wire dummy181;
SPLITT SplitCLK_4_1228(net1520,net1058_c1,dummy181);
wire dummy182;
SPLITT SplitCLK_2_1229(net1645,net1057_c1,dummy182);
wire dummy183;
SPLITT SplitCLK_2_1230(net1462,net1056_c1,dummy183);
wire dummy184;
SPLITT SplitCLK_2_1231(net2180,net1055_c1,dummy184);
wire dummy185;
SPLITT SplitCLK_2_1232(net2267,net1054_c1,dummy185);
wire dummy186;
SPLITT SplitCLK_4_1233(net1496,net1053_c1,dummy186);
wire dummy187;
SPLITT SplitCLK_2_1234(net2083,net1052_c1,dummy187);
wire dummy188;
SPLITT SplitCLK_2_1235(net2052,net1051_c1,dummy188);
wire dummy189;
SPLITT SplitCLK_2_1236(net1528,net1050_c1,dummy189);
wire dummy190;
SPLITT SplitCLK_2_1237(net2057,net1049_c1,dummy190);
wire dummy191;
SPLITT SplitCLK_2_1238(net1790,net1048_c1,dummy191);
wire dummy192;
SPLITT SplitCLK_4_1239(net2181,net1047_c1,dummy192);
wire dummy193;
SPLITT SplitCLK_4_1240(net2245,net1046_c1,dummy193);
wire dummy194;
SPLITT SplitCLK_2_1241(net1883,net1045_c1,dummy194);
wire dummy195;
SPLITT SplitCLK_2_1242(net2015,net1044_c1,dummy195);
wire dummy196;
SPLITT SplitCLK_2_1243(net1466,net1043_c1,dummy196);
wire dummy197;
SPLITT SplitCLK_2_1244(net1662,net1042_c1,dummy197);
wire dummy198;
SPLITT SplitCLK_4_1245(net1854,net1041_c1,dummy198);
wire dummy199;
SPLITT SplitCLK_4_1246(net1522,net1040_c1,dummy199);
wire dummy200;
SPLITT SplitCLK_2_1247(net1721,net1039_c1,dummy200);
wire dummy201;
SPLITT SplitCLK_4_1248(net1452,net1038_c1,dummy201);
wire dummy202;
SPLITT SplitCLK_2_1249(net1642,net1037_c1,dummy202);
wire dummy203;
SPLITT SplitCLK_2_1250(net2053,net1036_c1,dummy203);
wire dummy204;
SPLITT SplitCLK_2_1251(net1446,net1035_c1,dummy204);
wire dummy205;
SPLITT SplitCLK_2_1252(net1429,net1034_c1,dummy205);
wire dummy206;
SPLITT SplitCLK_2_1253(net1497,net1033_c1,dummy206);
wire dummy207;
SPLITT SplitCLK_4_1254(net1330,net1032_c1,dummy207);
wire dummy208;
SPLITT SplitCLK_2_1255(net1840,net1031_c1,dummy208);
wire dummy209;
SPLITT SplitCLK_2_1256(net1324,net1030_c1,dummy209);
wire dummy210;
SPLITT SplitCLK_4_1257(net1353,net1029_c1,dummy210);
wire dummy211;
SPLITT SplitCLK_2_1258(net1498,net1028_c1,dummy211);
wire dummy212;
SPLITT SplitCLK_2_1259(net1304,net1027_c1,dummy212);
wire dummy213;
SPLITT SplitCLK_2_1260(net1405,net1026_c1,dummy213);
wire dummy214;
SPLITT SplitCLK_2_1261(net1798,net1025_c1,dummy214);
wire dummy215;
SPLITT SplitCLK_2_1262(net1859,net1024_c1,dummy215);
wire dummy216;
SPLITT SplitCLK_2_1263(net1544,net1023_c1,dummy216);
wire dummy217;
SPLITT SplitCLK_2_1264(net1814,net1022_c1,dummy217);
wire dummy218;
SPLITT SplitCLK_4_1265(net1643,net1021_c1,dummy218);
wire dummy219;
SPLITT SplitCLK_4_1266(net1360,net1020_c1,dummy219);
wire dummy220;
SPLITT SplitCLK_2_1267(net1559,net1019_c1,dummy220);
wire dummy221;
SPLITT SplitCLK_4_1268(net1924,net1018_c1,dummy221);
wire dummy222;
SPLITT SplitCLK_2_1269(net2086,net1017_c1,dummy222);
wire dummy223;
SPLITT SplitCLK_2_1270(net1368,net1016_c1,dummy223);
wire dummy224;
SPLITT SplitCLK_2_1271(net1362,net1015_c1,dummy224);
wire dummy225;
SPLITT SplitCLK_2_1272(net1578,net1014_c1,dummy225);
wire dummy226;
SPLITT SplitCLK_4_1273(net1433,net1013_c1,dummy226);
wire dummy227;
SPLITT SplitCLK_4_1274(net1815,net1012_c1,dummy227);
wire dummy228;
SPLITT SplitCLK_2_1275(net1648,net1011_c1,dummy228);
wire dummy229;
SPLITT SplitCLK_4_1276(net1338,net1010_c1,dummy229);
wire dummy230;
SPLITT SplitCLK_2_1277(net1547,net1009_c1,dummy230);
wire dummy231;
SPLITT SplitCLK_2_1278(net1936,net1008_c1,dummy231);
wire dummy232;
SPLITT SplitCLK_4_1279(net2081,net1007_c1,dummy232);
wire dummy233;
SPLITT SplitCLK_2_1280(net1367,net1006_c1,dummy233);
wire dummy234;
SPLITT SplitCLK_4_1281(net1363,net1005_c1,dummy234);
wire dummy235;
SPLITT SplitCLK_4_1282(net1579,net1004_c1,dummy235);
wire dummy236;
SPLITT SplitCLK_4_1283(net2112,net1003_c1,dummy236);
wire dummy237;
SPLITT SplitCLK_2_1284(net1421,net1002_c1,dummy237);
wire dummy238;
SPLITT SplitCLK_2_1285(net1906,net1001_c1,dummy238);
wire dummy239;
SPLITT SplitCLK_2_1286(net1468,net1000_c1,dummy239);
wire dummy240;
SPLITT SplitCLK_2_1287(net1461,net999_c1,dummy240);
wire dummy241;
SPLITT SplitCLK_2_1288(net1553,net998_c1,dummy241);
wire dummy242;
SPLITT SplitCLK_4_1289(net1467,net997_c1,dummy242);
wire dummy243;
SPLITT SplitCLK_4_1290(net1514,net996_c1,dummy243);
wire dummy244;
SPLITT SplitCLK_4_1291(net1948,net995_c1,dummy244);
wire dummy245;
SPLITT SplitCLK_4_1292(net2194,net994_c1,dummy245);
wire dummy246;
SPLITT SplitCLK_2_1293(net2068,net993_c1,dummy246);
wire dummy247;
SPLITT SplitCLK_2_1294(net1884,net992_c1,dummy247);
wire dummy248;
SPLITT SplitCLK_4_1295(net1545,net991_c1,dummy248);
wire dummy249;
SPLITT SplitCLK_4_1296(net1612,net990_c1,dummy249);
wire dummy250;
SPLITT SplitCLK_2_1297(net2236,net989_c1,dummy250);
wire dummy251;
SPLITT SplitCLK_2_1298(net2118,net988_c1,dummy251);
wire dummy252;
SPLITT SplitCLK_2_1299(net1298,net987_c1,dummy252);
wire dummy253;
SPLITT SplitCLK_2_1300(net1415,net986_c1,dummy253);
wire dummy254;
SPLITT SplitCLK_4_1301(net1907,net985_c1,dummy254);
wire dummy255;
SPLITT SplitCLK_4_1302(net1649,net984_c1,dummy255);
wire dummy256;
SPLITT SplitCLK_4_1303(net1529,net983_c1,dummy256);
wire dummy257;
SPLITT SplitCLK_2_1304(net1339,net982_c1,dummy257);
wire dummy258;
SPLITT SplitCLK_4_1305(net1927,net981_c1,dummy258);
wire dummy259;
SPLITT SplitCLK_2_1306(net2020,net980_c1,dummy259);
wire dummy260;
SPLITT SplitCLK_4_1307(net2210,net979_c1,dummy260);
wire dummy261;
SPLITT SplitCLK_4_1308(net1885,net978_c1,dummy261);
wire dummy262;
SPLITT SplitCLK_2_1309(net1337,net977_c1,dummy262);
wire dummy263;
SPLITT SplitCLK_2_1310(net1707,net976_c1,dummy263);
wire dummy264;
SPLITT SplitCLK_4_1311(net2230,net975_c1,dummy264);
wire dummy265;
SPLITT SplitCLK_2_1312(net2243,net974_c1,dummy265);
wire dummy266;
SPLITT SplitCLK_4_1313(net1274,net973_c1,dummy266);
wire dummy267;
SPLITT SplitCLK_2_1314(net1427,net972_c1,dummy267);
wire dummy268;
SPLITT SplitCLK_2_1315(net1912,net971_c1,dummy268);
wire dummy269;
SPLITT SplitCLK_4_1316(net1463,net970_c1,dummy269);
wire dummy270;
SPLITT SplitCLK_2_1317(net1535,net969_c1,dummy270);
wire dummy271;
SPLITT SplitCLK_2_1318(net1270,net968_c1,dummy271);
wire dummy272;
SPLITT SplitCLK_2_1319(net2166,net967_c1,dummy272);
wire dummy273;
SPLITT SplitCLK_2_1320(net1332,net966_c1,dummy273);
wire dummy274;
SPLITT SplitCLK_2_1321(net1949,net965_c1,dummy274);
wire dummy275;
SPLITT SplitCLK_2_1322(net2164,net964_c1,dummy275);
wire dummy276;
SPLITT SplitCLK_2_1323(net1418,net963_c1,dummy276);
wire dummy277;
SPLITT SplitCLK_2_1324(net2208,net962_c1,dummy277);
wire dummy278;
SPLITT SplitCLK_4_1325(net1361,net961_c1,dummy278);
wire dummy279;
SPLITT SplitCLK_4_1326(net2273,net960_c1,dummy279);
wire dummy280;
SPLITT SplitCLK_4_1327(net1606,net959_c1,dummy280);
wire dummy281;
SPLITT SplitCLK_2_1328(net2231,net958_c1,dummy281);
wire dummy282;
SPLITT SplitCLK_2_1329(net2249,net957_c1,dummy282);
wire dummy283;
SPLITT SplitCLK_4_1330(net1584,net956_c1,dummy283);
wire dummy284;
SPLITT SplitCLK_2_1331(net1413,net955_c1,dummy284);
wire dummy285;
SPLITT SplitCLK_4_1332(net1277,net954_c1,dummy285);
wire dummy286;
SPLITT SplitCLK_4_1333(net1402,net953_c1,dummy286);
wire dummy287;
SPLITT SplitCLK_4_1334(net1937,net952_c1,dummy287);
wire dummy288;
SPLITT SplitCLK_4_1335(net1448,net951_c1,dummy288);
wire dummy289;
SPLITT SplitCLK_2_1336(net1974,net950_c1,dummy289);
wire dummy290;
SPLITT SplitCLK_2_1337(net2074,net949_c1,dummy290);
wire dummy291;
SPLITT SplitCLK_4_1338(net1333,net948_c1,dummy291);
wire dummy292;
SPLITT SplitCLK_2_1339(net1523,net947_c1,dummy292);
wire dummy293;
SPLITT SplitCLK_4_1340(net2075,net946_c1,dummy293);
wire dummy294;
SPLITT SplitCLK_4_1341(net1419,net945_c1,dummy294);
wire dummy295;
SPLITT SplitCLK_2_1342(net2214,net944_c1,dummy295);
wire dummy296;
SPLITT SplitCLK_2_1343(net1985,net943_c1,dummy296);
wire dummy297;
SPLITT SplitCLK_2_1344(net1861,net942_c1,dummy297);
wire dummy298;
SPLITT SplitCLK_2_1345(net1674,net941_c1,dummy298);
wire dummy299;
SPLITT SplitCLK_2_1346(net1609,net940_c1,dummy299);
wire dummy300;
SPLITT SplitCLK_4_1347(net2137,net939_c1,dummy300);
wire dummy301;
SPLITT SplitCLK_2_1348(net2274,net938_c1,dummy301);
wire dummy302;
SPLITT SplitCLK_4_1349(net1713,net937_c1,dummy302);
wire dummy303;
SPLITT SplitCLK_4_1350(net1389,net936_c1,dummy303);
wire dummy304;
SPLITT SplitCLK_4_1351(net1271,net935_c1,dummy304);
wire dummy305;
SPLITT SplitCLK_2_1352(net1403,net934_c1,dummy305);
wire dummy306;
SPLITT SplitCLK_4_1353(net1913,net933_c1,dummy306);
wire dummy307;
SPLITT SplitCLK_2_1354(net1453,net932_c1,dummy307);
wire dummy308;
SPLITT SplitCLK_4_1355(net1853,net931_c1,dummy308);
wire dummy309;
SPLITT SplitCLK_4_1356(net1975,net930_c1,dummy309);
wire dummy310;
SPLITT SplitCLK_2_1357(net2038,net929_c1,dummy310);
wire dummy311;
SPLITT SplitCLK_4_1358(net2069,net928_c1,dummy311);
wire dummy312;
SPLITT SplitCLK_2_1359(net1331,net927_c1,dummy312);
wire dummy313;
SPLITT SplitCLK_2_1360(net1516,net926_c1,dummy313);
wire dummy314;
SPLITT SplitCLK_4_1361(net1876,net925_c1,dummy314);
wire dummy315;
SPLITT SplitCLK_2_1362(net2073,net924_c1,dummy315);
wire dummy316;
SPLITT SplitCLK_4_1363(net2167,net923_c1,dummy316);
wire dummy317;
SPLITT SplitCLK_2_1364(net2197,net922_c1,dummy317);
wire dummy318;
SPLITT SplitCLK_2_1365(net2211,net921_c1,dummy318);
wire dummy319;
SPLITT SplitCLK_4_1366(net2279,net920_c1,dummy319);
wire dummy320;
SPLITT SplitCLK_4_1367(net1675,net919_c1,dummy320);
wire dummy321;
SPLITT SplitCLK_2_1368(net1613,net918_c1,dummy321);
wire dummy322;
SPLITT SplitCLK_4_1369(net2229,net917_c1,dummy322);
wire dummy323;
SPLITT SplitCLK_4_1370(net1596,net916_c1,dummy323);
wire dummy324;
SPLITT SplitCLK_4_1371(net1255,net915_c1,dummy324);
wire dummy325;
SPLITT SplitCLK_4_1372(net1382,net914_c1,dummy325);
wire dummy326;
SPLITT SplitCLK_2_1373(net1301,net913_c1,dummy326);
wire dummy327;
SPLITT SplitCLK_4_1374(net1396,net912_c1,dummy327);
wire dummy328;
SPLITT SplitCLK_2_1375(net1925,net911_c1,dummy328);
wire dummy329;
SPLITT SplitCLK_4_1376(net2258,net910_c1,dummy329);
wire dummy330;
SPLITT SplitCLK_4_1377(net1888,net909_c1,dummy330);
wire dummy331;
SPLITT SplitCLK_4_1378(net1998,net908_c1,dummy331);
wire dummy332;
SPLITT SplitCLK_4_1379(net1673,net907_c1,dummy332);
wire dummy333;
SPLITT SplitCLK_2_1380(net2066,net906_c1,dummy333);
wire dummy334;
SPLITT SplitCLK_2_1381(net2186,net905_c1,dummy334);
wire dummy335;
SPLITT SplitCLK_2_1382(net1521,net904_c1,dummy335);
wire dummy336;
SPLITT SplitCLK_2_1383(net1874,net903_c1,dummy336);
wire dummy337;
SPLITT SplitCLK_2_1384(net1889,net902_c1,dummy337);
wire dummy338;
SPLITT SplitCLK_2_1385(net2172,net901_c1,dummy338);
wire dummy339;
SPLITT SplitCLK_4_1386(net2209,net900_c1,dummy339);
wire dummy340;
SPLITT SplitCLK_4_1387(net2087,net899_c1,dummy340);
wire dummy341;
SPLITT SplitCLK_4_1388(net2275,net898_c1,dummy341);
wire dummy342;
SPLITT SplitCLK_2_1389(net1680,net897_c1,dummy342);
wire dummy343;
SPLITT SplitCLK_4_1390(net1750,net896_c1,dummy343);
wire dummy344;
SPLITT SplitCLK_2_1391(net1709,net895_c1,dummy344);
wire dummy345;
SPLITT SplitCLK_4_1392(net1590,net894_c1,dummy345);
wire dummy346;
SPLITT SplitCLK_2_1393(net1383,net893_c1,dummy346);
wire dummy347;
SPLITT SplitCLK_2_1394(net1319,net892_c1,dummy347);
wire dummy348;
SPLITT SplitCLK_2_1395(net1397,net891_c1,dummy348);
wire dummy349;
SPLITT SplitCLK_4_1396(net1919,net890_c1,dummy349);
wire dummy350;
SPLITT SplitCLK_4_1397(net1560,net889_c1,dummy350);
wire dummy351;
SPLITT SplitCLK_2_1398(net1585,net888_c1,dummy351);
wire dummy352;
SPLITT SplitCLK_2_1399(net1622,net887_c1,dummy352);
wire dummy353;
SPLITT SplitCLK_4_1400(net2019,net886_c1,dummy353);
wire dummy354;
SPLITT SplitCLK_4_1401(net1877,net885_c1,dummy354);
wire dummy355;
SPLITT SplitCLK_4_1402(net1950,net884_c1,dummy355);
wire dummy356;
SPLITT SplitCLK_2_1403(net1844,net883_c1,dummy356);
wire dummy357;
SPLITT SplitCLK_2_1404(net1493,net882_c1,dummy357);
wire dummy358;
SPLITT SplitCLK_2_1405(net2067,net881_c1,dummy358);
wire dummy359;
SPLITT SplitCLK_4_1406(net2187,net880_c1,dummy359);
wire dummy360;
SPLITT SplitCLK_4_1407(net1517,net879_c1,dummy360);
wire dummy361;
SPLITT SplitCLK_4_1408(net1576,net878_c1,dummy361);
wire dummy362;
SPLITT SplitCLK_4_1409(net1871,net877_c1,dummy362);
wire dummy363;
SPLITT SplitCLK_4_1410(net1868,net876_c1,dummy363);
wire dummy364;
SPLITT SplitCLK_4_1411(net2173,net875_c1,dummy364);
wire dummy365;
SPLITT SplitCLK_4_1412(net2170,net874_c1,dummy365);
wire dummy366;
SPLITT SplitCLK_4_1413(net1681,net873_c1,dummy366);
wire dummy367;
SPLITT SplitCLK_2_1414(net1751,net872_c1,dummy367);
wire dummy368;
SPLITT SplitCLK_4_1415(net1566,net871_c1,dummy368);
wire dummy369;
SPLITT SplitCLK_2_1416(net1627,net870_c1,dummy369);
wire dummy370;
SPLITT SplitCLK_4_1417(net1290,net869_c1,dummy370);
wire dummy371;
SPLITT SplitCLK_2_1418(net1316,net868_c1,dummy371);
wire dummy372;
SPLITT SplitCLK_4_1419(net1305,net867_c1,dummy372);
wire dummy373;
SPLITT SplitCLK_4_1420(net2119,net866_c1,dummy373);
wire dummy374;
SPLITT SplitCLK_2_1421(net2113,net865_c1,dummy374);
wire dummy375;
SPLITT SplitCLK_2_1422(net1628,net864_c1,dummy375);
wire dummy376;
SPLITT SplitCLK_2_1423(net1776,net863_c1,dummy376);
wire dummy377;
SPLITT SplitCLK_2_1424(net1970,net862_c1,dummy377);
wire dummy378;
SPLITT SplitCLK_2_1425(net1951,net861_c1,dummy378);
wire dummy379;
SPLITT SplitCLK_4_1426(net1846,net860_c1,dummy379);
wire dummy380;
SPLITT SplitCLK_4_1427(net2042,net859_c1,dummy380);
wire dummy381;
SPLITT SplitCLK_2_1428(net2184,net858_c1,dummy381);
wire dummy382;
SPLITT SplitCLK_2_1429(net1515,net857_c1,dummy382);
wire dummy383;
SPLITT SplitCLK_4_1430(net1583,net856_c1,dummy383);
wire dummy384;
SPLITT SplitCLK_2_1431(net1890,net855_c1,dummy384);
wire dummy385;
SPLITT SplitCLK_4_1432(net1875,net854_c1,dummy385);
wire dummy386;
SPLITT SplitCLK_4_1433(net2185,net853_c1,dummy386);
wire dummy387;
SPLITT SplitCLK_2_1434(net2195,net852_c1,dummy387);
wire dummy388;
SPLITT SplitCLK_4_1435(net1757,net851_c1,dummy388);
wire dummy389;
SPLITT SplitCLK_2_1436(net2051,net850_c1,dummy389);
wire dummy390;
SPLITT SplitCLK_2_1437(net1727,net849_c1,dummy390);
wire dummy391;
SPLITT SplitCLK_2_1438(net1567,net848_c1,dummy391);
wire dummy392;
SPLITT SplitCLK_4_1439(net1623,net847_c1,dummy392);
wire dummy393;
SPLITT SplitCLK_2_1440(net1291,net846_c1,dummy393);
wire dummy394;
SPLITT SplitCLK_4_1441(net1317,net845_c1,dummy394);
wire dummy395;
SPLITT SplitCLK_4_1442(net1299,net844_c1,dummy395);
wire dummy396;
SPLITT SplitCLK_2_1443(net2142,net843_c1,dummy396);
wire dummy397;
SPLITT SplitCLK_4_1444(net1905,net842_c1,dummy397);
wire dummy398;
SPLITT SplitCLK_4_1445(net1777,net841_c1,dummy398);
wire dummy399;
SPLITT SplitCLK_2_1446(net1983,net840_c1,dummy399);
wire dummy400;
SPLITT SplitCLK_4_1447(net2001,net839_c1,dummy400);
wire dummy401;
SPLITT SplitCLK_4_1448(net1384,net838_c1,dummy401);
wire dummy402;
SPLITT SplitCLK_2_1449(net1869,net837_c1,dummy402);
wire dummy403;
SPLITT SplitCLK_2_1450(net2036,net836_c1,dummy403);
wire dummy404;
SPLITT SplitCLK_4_1451(net1663,net835_c1,dummy404);
wire dummy405;
SPLITT SplitCLK_4_1452(net2178,net834_c1,dummy405);
wire dummy406;
SPLITT SplitCLK_2_1453(net1828,net833_c1,dummy406);
wire dummy407;
SPLITT SplitCLK_2_1454(net1561,net832_c1,dummy407);
wire dummy408;
SPLITT SplitCLK_2_1455(net1455,net831_c1,dummy408);
wire dummy409;
SPLITT SplitCLK_2_1456(net1829,net830_c1,dummy409);
wire dummy410;
SPLITT SplitCLK_2_1457(net2171,net829_c1,dummy410);
wire dummy411;
SPLITT SplitCLK_2_1458(net1745,net828_c1,dummy411);
wire dummy412;
SPLITT SplitCLK_4_1459(net2105,net827_c1,dummy412);
wire dummy413;
SPLITT SplitCLK_2_1460(net2131,net826_c1,dummy413);
wire dummy414;
SPLITT SplitCLK_2_1461(net1597,net825_c1,dummy414);
wire dummy415;
SPLITT SplitCLK_4_1462(net1286,net824_c1,dummy415);
wire dummy416;
SPLITT SplitCLK_2_1463(net1323,net823_c1,dummy416);
wire dummy417;
SPLITT SplitCLK_2_1464(net1399,net822_c1,dummy417);
wire dummy418;
SPLITT SplitCLK_4_1465(net1845,net821_c1,dummy418);
wire dummy419;
SPLITT SplitCLK_4_1466(net1355,net820_c1,dummy419);
wire dummy420;
SPLITT SplitCLK_2_1467(net2045,net819_c1,dummy420);
wire dummy421;
SPLITT SplitCLK_2_1468(net1659,net818_c1,dummy421);
wire dummy422;
SPLITT SplitCLK_2_1469(net1621,net817_c1,dummy422);
wire dummy423;
SPLITT SplitCLK_4_1470(net2143,net816_c1,dummy423);
wire dummy424;
SPLITT SplitCLK_4_1471(net2235,net815_c1,dummy424);
wire dummy425;
SPLITT SplitCLK_4_1472(net1752,net814_c1,dummy425);
wire dummy426;
SPLITT SplitCLK_2_1473(net2114,net813_c1,dummy426);
wire dummy427;
SPLITT SplitCLK_2_1474(net1910,net812_c1,dummy427);
wire dummy428;
SPLITT SplitCLK_2_1475(net1782,net811_c1,dummy428);
wire dummy429;
SPLITT SplitCLK_2_1476(net1989,net810_c1,dummy429);
wire dummy430;
SPLITT SplitCLK_2_1477(net1999,net809_c1,dummy430);
wire dummy431;
SPLITT SplitCLK_2_1478(net1385,net808_c1,dummy431);
wire dummy432;
SPLITT SplitCLK_2_1479(net1847,net807_c1,dummy432);
wire dummy433;
SPLITT SplitCLK_4_1480(net2037,net806_c1,dummy433);
wire dummy434;
SPLITT SplitCLK_2_1481(net1678,net805_c1,dummy434);
wire dummy435;
SPLITT SplitCLK_2_1482(net2179,net804_c1,dummy435);
wire dummy436;
SPLITT SplitCLK_4_1483(net1822,net803_c1,dummy436);
wire dummy437;
SPLITT SplitCLK_2_1484(net1607,net802_c1,dummy437);
wire dummy438;
SPLITT SplitCLK_2_1485(net1449,net801_c1,dummy438);
wire dummy439;
SPLITT SplitCLK_4_1486(net1968,net800_c1,dummy439);
wire dummy440;
SPLITT SplitCLK_4_1487(net2165,net799_c1,dummy440);
wire dummy441;
SPLITT SplitCLK_2_1488(net2101,net798_c1,dummy441);
wire dummy442;
SPLITT SplitCLK_2_1489(net2280,net797_c1,dummy442);
wire dummy443;
SPLITT SplitCLK_2_1490(net2260,net796_c1,dummy443);
wire dummy444;
SPLITT SplitCLK_4_1491(net1592,net795_c1,dummy444);
wire dummy445;
SPLITT SplitCLK_4_1492(net1284,net794_c1,dummy445);
wire dummy446;
SPLITT SplitCLK_4_1493(net1325,net793_c1,dummy446);
wire dummy447;
SPLITT SplitCLK_2_1494(net1753,net792_c1,dummy447);
wire dummy448;
SPLITT SplitCLK_4_1495(net2115,net791_c1,dummy448);
wire dummy449;
SPLITT SplitCLK_2_1496(net2216,net790_c1,dummy449);
wire dummy450;
SPLITT SplitCLK_4_1497(net1911,net789_c1,dummy450);
wire dummy451;
SPLITT SplitCLK_4_1498(net1783,net788_c1,dummy451);
wire dummy452;
SPLITT SplitCLK_4_1499(net1991,net787_c1,dummy452);
wire dummy453;
SPLITT SplitCLK_4_1500(net1976,net786_c1,dummy453);
wire dummy454;
SPLITT SplitCLK_4_1501(net1268,net785_c1,dummy454);
wire dummy455;
SPLITT SplitCLK_4_1502(net1292,net784_c1,dummy455);
wire dummy456;
SPLITT SplitCLK_4_1503(net1841,net783_c1,dummy456);
wire dummy457;
SPLITT SplitCLK_2_1504(net2043,net782_c1,dummy457);
wire dummy458;
SPLITT SplitCLK_4_1505(net1679,net781_c1,dummy458);
wire dummy459;
SPLITT SplitCLK_2_1506(net1823,net780_c1,dummy459);
wire dummy460;
SPLITT SplitCLK_2_1507(net1577,net779_c1,dummy460);
wire dummy461;
SPLITT SplitCLK_4_1508(net1447,net778_c1,dummy461);
wire dummy462;
SPLITT SplitCLK_4_1509(net1971,net777_c1,dummy462);
wire dummy463;
SPLITT SplitCLK_4_1510(net2237,net776_c1,dummy463);
wire dummy464;
SPLITT SplitCLK_2_1511(net1591,net775_c1,dummy464);
wire dummy465;
SPLITT SplitCLK_2_1512(net1285,net774_c1,dummy465);
wire dummy466;
SPLITT SplitCLK_4_1513(net1728,net773_c1,dummy466);
wire dummy467;
SPLITT SplitCLK_2_1514(net2120,net772_c1,dummy467);
wire dummy468;
SPLITT SplitCLK_2_1515(net1934,net771_c1,dummy468);
wire dummy469;
SPLITT SplitCLK_2_1516(net1806,net770_c1,dummy469);
wire dummy470;
SPLITT SplitCLK_2_1517(net2013,net769_c1,dummy470);
wire dummy471;
SPLITT SplitCLK_2_1518(net1977,net768_c1,dummy471);
wire dummy472;
SPLITT SplitCLK_2_1519(net1275,net767_c1,dummy472);
wire dummy473;
SPLITT SplitCLK_2_1520(net1293,net766_c1,dummy473);
wire dummy474;
SPLITT SplitCLK_2_1521(net1484,net765_c1,dummy474);
wire dummy475;
SPLITT SplitCLK_4_1522(net1469,net764_c1,dummy475);
wire dummy476;
SPLITT SplitCLK_4_1523(net2039,net763_c1,dummy476);
wire dummy477;
SPLITT SplitCLK_4_1524(net1799,net762_c1,dummy477);
wire dummy478;
SPLITT SplitCLK_4_1525(net1737,net761_c1,dummy478);
wire dummy479;
SPLITT SplitCLK_2_1526(net1743,net760_c1,dummy479);
wire dummy480;
SPLITT SplitCLK_2_1527(net1969,net759_c1,dummy480);
wire dummy481;
SPLITT SplitCLK_2_1528(net2259,net758_c1,dummy481);
wire dummy482;
SPLITT SplitCLK_2_1529(net1593,net757_c1,dummy482);
wire dummy483;
SPLITT SplitCLK_4_1530(net1261,net756_c1,dummy483);
wire dummy484;
SPLITT SplitCLK_2_1531(net1729,net755_c1,dummy484);
wire dummy485;
SPLITT SplitCLK_4_1532(net2121,net754_c1,dummy485);
wire dummy486;
SPLITT SplitCLK_4_1533(net2215,net753_c1,dummy486);
wire dummy487;
SPLITT SplitCLK_4_1534(net1935,net752_c1,dummy487);
wire dummy488;
SPLITT SplitCLK_4_1535(net1807,net751_c1,dummy488);
wire dummy489;
SPLITT SplitCLK_2_1536(net2007,net750_c1,dummy489);
wire dummy490;
SPLITT SplitCLK_2_1537(net1434,net749_c1,dummy490);
wire dummy491;
SPLITT SplitCLK_2_1538(net1269,net748_c1,dummy491);
wire dummy492;
SPLITT SplitCLK_2_1539(net1287,net747_c1,dummy492);
wire dummy493;
SPLITT SplitCLK_4_1540(net1485,net746_c1,dummy493);
wire dummy494;
SPLITT SplitCLK_2_1541(net1855,net745_c1,dummy494);
wire dummy495;
SPLITT SplitCLK_2_1542(net2059,net744_c1,dummy495);
wire dummy496;
SPLITT SplitCLK_4_1543(net1791,net743_c1,dummy496);
wire dummy497;
SPLITT SplitCLK_4_1544(net1531,net742_c1,dummy497);
wire dummy498;
SPLITT SplitCLK_2_1545(net2261,net741_c1,dummy498);
wire dummy499;
SPLITT SplitCLK_2_1546(net1599,net740_c1,dummy499);
SPLITT SplitCLK_0_1547(net2284,net738_c1,net739_c1);
wire dummy500;
SPLITT Split_HOLD_1667(net553,dummy500,net2285_c1);
wire dummy501;
SPLITT Split_HOLD_1668(net496,dummy501,net2286_c1);
wire dummy502;
SPLITT Split_HOLD_1669(net490,dummy502,net2287_c1);
wire dummy503;
SPLITT Split_HOLD_1670(net484,dummy503,net2288_c1);
wire dummy504;
SPLITT Split_HOLD_1671(net712,dummy504,net2289_c1);
wire dummy505;
SPLITT Split_HOLD_1672(net454,dummy505,net2290_c1);
wire dummy506;
SPLITT Split_HOLD_1673(net411,dummy506,net2291_c1);
wire dummy507;
SPLITT Split_HOLD_1674(net667,dummy507,net2292_c1);
wire dummy508;
SPLITT Split_HOLD_1675(net658,dummy508,net2293_c1);
wire dummy509;
SPLITT Split_HOLD_1676(net363,dummy509,net2294_c1);
wire dummy510;
SPLITT Split_HOLD_1677(net633,dummy510,net2295_c1);
wire dummy511;
SPLITT Split_HOLD_1678(net353,dummy511,net2296_c1);
wire dummy512;
SPLITT Split_HOLD_1679(net597,dummy512,net2297_c1);
wire dummy513;
SPLITT Split_HOLD_1680(net685,dummy513,net2298_c1);
wire dummy514;
SPLITT Split_HOLD_1681(net660,dummy514,net2299_c1);
wire dummy515;
SPLITT Split_HOLD_1682(net631,dummy515,net2300_c1);
wire dummy516;
SPLITT Split_HOLD_1683(net610,dummy516,net2301_c1);
wire dummy517;
SPLITT Split_HOLD_1684(net607,dummy517,net2302_c1);
wire dummy518;
SPLITT Split_HOLD_1685(net347,dummy518,net2303_c1);
INTERCONNECT D0_Pad_Split_552_n1732(D0_Pad,net0);
INTERCONNECT D1_Pad_Split_549_n1729(D1_Pad,net1);
INTERCONNECT D2_Pad_Split_548_n1728(D2_Pad,net2);
INTERCONNECT D3_Pad_Split_546_n1726(D3_Pad,net3);
INTERCONNECT DFFT_540_Q0_Q0_Pad(net4_c1,Q0_Pad);
INTERCONNECT DFFT_538_Q1_Q1_Pad(net5_c1,Q1_Pad);
INTERCONNECT XOR2T_134_R0_R0_Pad(net6_c1,R0_Pad);
INTERCONNECT DFFT_527_Q2_Q2_Pad(net7_c1,Q2_Pad);
INTERCONNECT OR2T_133_R1_R1_Pad(net8_c1,R1_Pad);
INTERCONNECT DFFT_511_Q3_Q3_Pad(net9_c1,Q3_Pad);
INTERCONNECT OR2T_127_R2_R2_Pad(net10_c1,R2_Pad);
INTERCONNECT AND2T_120_R3_R3_Pad(net11_c1,R3_Pad);
INTERCONNECT X0_Pad_Split_545_n1725(X0_Pad,net12);
INTERCONNECT X1_Pad_Split_543_n1723(X1_Pad,net13);
INTERCONNECT X2_Pad_Split_542_n1722(X2_Pad,net14);
INTERCONNECT X3_Pad_Split_541_n1721(X3_Pad,net15);
INTERCONNECT NOTT_20_n20_Split_558_n1738(net16_c1,net16);
INTERCONNECT NOTT_21_n21_OR2T_80_n81(net17_c1,net17);
INTERCONNECT AND2T_29_n30_Split_562_n1742(net18_c1,net18);
INTERCONNECT OR2T_22_n22_AND2T_23_n23(net19_c1,net19);
INTERCONNECT OR2T_30_n31_AND2T_29_n30(net20_c1,net20);
INTERCONNECT AND2T_23_n23_AND2T_24_n24(net21_c1,net21);
INTERCONNECT OR2T_39_n40_DFFT_162__FPB_n1342(net22_c1,net22);
INTERCONNECT OR2T_31_n32_OR2T_34_n35(net23_c1,net23);
INTERCONNECT AND2T_24_n24_DFFT_496__FPB_n1676(net24_c1,net24);
INTERCONNECT OR2T_40_n41_AND2T_43_n44(net25_c1,net25);
INTERCONNECT NOTT_32_n33_DFFT_294__FPB_n1474(net26_c1,net26);
INTERCONNECT OR2T_25_n25_Split_559_n1739(net27_c1,net27);
INTERCONNECT NOTT_17_n17_Split_554_n1734(net28_c1,net28);
INTERCONNECT AND2T_49_n50_AND2T_50_n51(net29_c1,net29);
INTERCONNECT OR2T_41_n42_AND2T_42_n43(net30_c1,net30);
INTERCONNECT AND2T_33_n34_OR2T_34_n35(net31_c1,net31);
INTERCONNECT OR2T_26_n26_AND2T_27_n27(net32_c1,net32);
INTERCONNECT NOTT_18_n18_DFFT_325__FPB_n1505(net33_c1,net33);
INTERCONNECT AND2T_50_n51_OR2T_51_n52(net34_c1,net34);
INTERCONNECT AND2T_42_n43_AND2T_43_n44(net35_c1,net35);
INTERCONNECT OR2T_34_n35_Split_564_n1744(net36_c1,net36);
INTERCONNECT AND2T_27_n27_Split_560_n1740(net37_c1,net37);
INTERCONNECT AND2T_19_n19_Split_556_n1736(net38_c1,net38);
INTERCONNECT AND2T_59_n60_OR2T_64_n65(net39_c1,net39);
INTERCONNECT OR2T_51_n52_OR2T_52_n53(net40_c1,net40);
INTERCONNECT AND2T_43_n44_Split_569_n1749(net41_c1,net41);
INTERCONNECT AND2T_35_n36_Split_566_n1746(net42_c1,net42);
INTERCONNECT AND2T_28_n28_Split_561_n1741(net43_c1,net43);
INTERCONNECT OR2T_60_n61_AND2T_59_n60(net44_c1,net44);
INTERCONNECT OR2T_52_n53_Split_571_n1751(net45_c1,net45);
INTERCONNECT XOR2T_44_n45_OR2T_51_n52(net46_c1,net46);
INTERCONNECT OR2T_36_n37_AND2T_35_n36(net47_c1,net47);
INTERCONNECT AND2T_69_n70_Split_584_n1764(net48_c1,net48);
INTERCONNECT AND2T_61_n62_OR2T_63_n64(net49_c1,net49);
INTERCONNECT AND2T_53_n54_Split_573_n1753(net50_c1,net50);
INTERCONNECT OR2T_45_n46_XOR2T_44_n45(net51_c1,net51);
INTERCONNECT OR2T_37_n38_Split_567_n1747(net52_c1,net52);
INTERCONNECT NOTT_70_n71_AND2T_69_n70(net53_c1,net53);
INTERCONNECT XOR2T_62_n63_DFFT_192__FPB_n1372(net54_c1,net54);
INTERCONNECT AND2T_54_n55_Split_575_n1755(net55_c1,net55);
INTERCONNECT OR2T_46_n47_AND2T_50_n51(net56_c1,net56);
INTERCONNECT AND2T_38_n39_Split_568_n1748(net57_c1,net57);
INTERCONNECT OR2T_79_n80_DFFT_273__FPB_n1453(net58_c1,net58);
INTERCONNECT OR2T_71_n72_Split_587_n1767(net59_c1,net59);
INTERCONNECT OR2T_63_n64_OR2T_64_n65(net60_c1,net60);
INTERCONNECT NOTT_55_n56_Split_576_n1756(net61_c1,net61);
INTERCONNECT XOR2T_47_n48_DFFT_178__FPB_n1358(net62_c1,net62);
INTERCONNECT OR2T_80_n81_Split_593_n1773(net63_c1,net63);
INTERCONNECT XOR2T_72_n73_Split_588_n1768(net64_c1,net64);
INTERCONNECT OR2T_64_n65_Split_582_n1762(net65_c1,net65);
INTERCONNECT NOTT_56_n57_Split_579_n1759(net66_c1,net66);
INTERCONNECT OR2T_48_n49_AND2T_49_n50(net67_c1,net67);
INTERCONNECT XOR2T_89_n90_XOR2T_91_n92(net68_c1,net68);
INTERCONNECT OR2T_81_n82_Split_595_n1775(net69_c1,net69);
INTERCONNECT OR2T_73_n74_Split_589_n1769(net70_c1,net70);
INTERCONNECT XOR2T_65_n66_DFFT_201__FPB_n1381(net71_c1,net71);
INTERCONNECT AND2T_57_n58_DFFT_196__FPB_n1376(net72_c1,net72);
INTERCONNECT OR2T_90_n91_XOR2T_89_n90(net73_c1,net73);
INTERCONNECT AND2T_82_n83_Split_596_n1776(net74_c1,net74);
INTERCONNECT XOR2T_74_n75_DFFT_238__FPB_n1418(net75_c1,net75);
INTERCONNECT AND2T_66_n67_XOR2T_65_n66(net76_c1,net76);
INTERCONNECT NOTT_58_n59_Split_581_n1761(net77_c1,net77);
INTERCONNECT XOR2T_91_n92_DFFT_285__FPB_n1465(net78_c1,net78);
INTERCONNECT NOTT_83_n84_AND2T_82_n83(net79_c1,net79);
INTERCONNECT AND2T_75_n76_DFFT_239__FPB_n1419(net80_c1,net80);
INTERCONNECT AND2T_67_n68_NOTT_70_n71(net81_c1,net81);
INTERCONNECT AND2T_92_n93_NOTT_94_n95(net82_c1,net82);
INTERCONNECT OR2T_84_n85_AND2T_85_n86(net83_c1,net83);
INTERCONNECT AND2T_76_n77_Split_590_n1770(net84_c1,net84);
INTERCONNECT OR2T_68_n69_DFFT_206__FPB_n1386(net85_c1,net85);
INTERCONNECT XOR2T_93_n94_AND2T_92_n93(net86_c1,net86);
INTERCONNECT AND2T_85_n86_OR2T_86_n87(net87_c1,net87);
INTERCONNECT NOTT_77_n78_AND2T_78_n79(net88_c1,net88);
INTERCONNECT NOTT_94_n95_Split_597_n1777(net89_c1,net89);
INTERCONNECT OR2T_86_n87_AND2T_87_n88(net90_c1,net90);
INTERCONNECT AND2T_78_n79_Split_592_n1772(net91_c1,net91);
INTERCONNECT AND2T_95_n96_XOR2T_100_n101(net92_c1,net92);
INTERCONNECT AND2T_87_n88_OR2T_102_n103(net93_c1,net93);
INTERCONNECT OR2T_96_n97_NOTT_97_n98(net94_c1,net94);
INTERCONNECT AND2T_88_n89_XOR2T_93_n94(net95_c1,net95);
INTERCONNECT NOTT_97_n98_DFFT_296__FPB_n1476(net96_c1,net96);
INTERCONNECT OR2T_98_n99_Split_598_n1778(net97_c1,net97);
INTERCONNECT AND2T_99_n100_DFFT_308__FPB_n1488(net98_c1,net98);
INTERCONNECT XOR2T_100_n101_Split_599_n1779(net99_c1,net99);
INTERCONNECT AND2T_109_n110_Split_603_n1783(net100_c1,net100);
INTERCONNECT NOTT_101_n102_DFFT_309__FPB_n1489(net101_c1,net101);
INTERCONNECT NOTT_110_n111_DFFT_359__FPB_n1539(net102_c1,net102);
INTERCONNECT OR2T_102_n103_Split_601_n1781(net103_c1,net103);
INTERCONNECT OR2T_119_n120_AND2T_120_R3(net104_c1,net104);
INTERCONNECT OR2T_111_n112_AND2T_112_n113(net105_c1,net105);
INTERCONNECT AND2T_103_n104_AND2T_135_n136(net106_c1,net106);
INTERCONNECT AND2T_112_n113_Split_604_n1784(net107_c1,net107);
INTERCONNECT NOTT_104_n105_DFFT_368__FPB_n1548(net108_c1,net108);
INTERCONNECT AND2T_129_n130_DFFT_430__FPB_n1610(net109_c1,net109);
INTERCONNECT NOTT_121_n122_AND2T_120_R3(net110_c1,net110);
INTERCONNECT OR2T_113_n114_Split_605_n1785(net111_c1,net111);
INTERCONNECT XOR2T_105_n106_DFFT_367__FPB_n1547(net112_c1,net112);
INTERCONNECT OR2T_130_n131_DFFT_431__FPB_n1611(net113_c1,net113);
INTERCONNECT XOR2T_122_n123_DFFT_394__FPB_n1574(net114_c1,net114);
INTERCONNECT AND2T_114_n115_OR2T_115_n116(net115_c1,net115);
INTERCONNECT AND2T_106_n107_Split_602_n1782(net116_c1,net116);
INTERCONNECT NOTT_139_n140_Split_617_n1797(net117_c1,net117);
INTERCONNECT AND2T_131_n132_OR2T_133_R1(net118_c1,net118);
INTERCONNECT AND2T_123_n124_OR2T_127_R2(net119_c1,net119);
INTERCONNECT OR2T_115_n116_Split_606_n1786(net120_c1,net120);
INTERCONNECT NOTT_107_n108_AND2T_106_n107(net121_c1,net121);
INTERCONNECT AND2T_140_n141_Split_620_n1800(net122_c1,net122);
INTERCONNECT AND2T_132_n133_OR2T_133_R1(net123_c1,net123);
INTERCONNECT AND2T_124_n125_OR2T_125_n126(net124_c1,net124);
INTERCONNECT AND2T_116_n117_NOTT_121_n122(net125_c1,net125);
INTERCONNECT OR2T_108_n109_AND2T_109_n110(net126_c1,net126);
INTERCONNECT AND2T_141_n142_Split_623_n1803(net127_c1,net127);
INTERCONNECT OR2T_125_n126_Split_607_n1787(net128_c1,net128);
INTERCONNECT XOR2T_117_n118_AND2T_116_n117(net129_c1,net129);
INTERCONNECT AND2T_126_n127_OR2T_127_R2(net130_c1,net130);
INTERCONNECT AND2T_118_n119_DFFT_387__FPB_n1567(net131_c1,net131);
INTERCONNECT AND2T_135_n136_XOR2T_134_R0(net132_c1,net132);
INTERCONNECT NOTT_136_n137_Split_608_n1788(net133_c1,net133);
INTERCONNECT XOR2T_128_n129_OR2T_130_n131(net134_c1,net134);
INTERCONNECT NOTT_137_n138_Split_611_n1791(net135_c1,net135);
INTERCONNECT NOTT_138_n139_Split_614_n1794(net136_c1,net136);
INTERCONNECT Split_620_n1800_Split_622_n1802(net137_c1,net137);
INTERCONNECT Split_541_n1721_DFFT_142__FPB_n143(net138_c1,net138);
INTERCONNECT Split_621_n1801_OR2T_68_n69(net139_c1,net139);
INTERCONNECT Split_550_n1730_DFFT_145__FPB_n146(net140_c1,net140);
INTERCONNECT Split_622_n1802_DFFT_528__FPB_n1708(net141_c1,net141);
INTERCONNECT Split_542_n1722_DFFT_143__FPB_n144(net142_c1,net142);
INTERCONNECT Split_630_n1810_XOR2T_47_n48(net143_c1,net143);
INTERCONNECT Split_623_n1803_Split_625_n1805(net144_c1,net144);
INTERCONNECT Split_551_n1731_DFFT_346__FPB_n1526(net145_c1,net145);
INTERCONNECT Split_543_n1723_Split_544_n1724(net146_c1,net146);
INTERCONNECT Split_631_n1811_DFFT_175__FPB_n1355(net147_c1,net147);
INTERCONNECT Split_632_n1812_Split_634_n1814(net148_c1,net148);
INTERCONNECT Split_552_n1732_Split_553_n1733(net149_c1,net149);
INTERCONNECT Split_624_n1804_AND2T_123_n124(net150_c1,net150);
INTERCONNECT Split_544_n1724_DFFT_166__FPB_n1346(net151_c1,net151);
INTERCONNECT Split_640_n1820_AND2T_57_n58(net152_c1,net152);
INTERCONNECT Split_560_n1740_AND2T_61_n62(net153_c1,net153);
INTERCONNECT Split_641_n1821_Split_643_n1823(net154_c1,net154);
INTERCONNECT Split_545_n1725_DFFT_441__FPB_n1621(net155_c1,net155);
INTERCONNECT Split_553_n1733_DFFT_146__FPB_n147(net156_c1,net156);
INTERCONNECT Split_625_n1805_DFFT_539__FPB_n1719(net157_c1,net157);
INTERCONNECT Split_561_n1741_DFFT_512__FPB_n1692(net158_c1,net158);
INTERCONNECT Split_633_n1813_OR2T_31_n32(net159_c1,net159);
INTERCONNECT Split_626_n1806_Split_628_n1808(net160_c1,net160);
INTERCONNECT Split_562_n1742_Split_563_n1743(net161_c1,net161);
INTERCONNECT Split_554_n1734_Split_555_n1735(net162_c1,net162);
INTERCONNECT Split_634_n1814_DFFT_278__FPB_n1458(net163_c1,net163);
INTERCONNECT Split_546_n1726_Split_547_n1727(net164_c1,net164);
INTERCONNECT Split_642_n1822_XOR2T_74_n75(net165_c1,net165);
INTERCONNECT Split_570_n1750_OR2T_90_n91(net166_c1,net166);
INTERCONNECT Split_635_n1815_Split_637_n1817(net167_c1,net167);
INTERCONNECT Split_643_n1823_DFFT_460__FPB_n1640(net168_c1,net168);
INTERCONNECT Split_571_n1751_Split_572_n1752(net169_c1,net169);
INTERCONNECT Split_563_n1743_DFFT_181__FPB_n1361(net170_c1,net170);
INTERCONNECT Split_627_n1807_OR2T_26_n26(net171_c1,net171);
INTERCONNECT Split_555_n1735_DFFT_151__FPB_n1331(net172_c1,net172);
INTERCONNECT Split_547_n1727_DFFT_152__FPB_n1332(net173_c1,net173);
INTERCONNECT Split_556_n1736_Split_557_n1737(net174_c1,net174);
INTERCONNECT Split_548_n1728_DFFT_144__FPB_n145(net175_c1,net175);
INTERCONNECT Split_564_n1744_Split_565_n1745(net176_c1,net176);
INTERCONNECT Split_580_n1760_XOR2T_74_n75(net177_c1,net177);
INTERCONNECT Split_572_n1752_AND2T_76_n77(net178_c1,net178);
INTERCONNECT Split_628_n1808_NOTT_32_n33(net179_c1,net179);
INTERCONNECT Split_636_n1816_AND2T_33_n34(net180_c1,net180);
INTERCONNECT Split_629_n1809_Split_631_n1811(net181_c1,net181);
INTERCONNECT Split_549_n1729_Split_551_n1731(net182_c1,net182);
INTERCONNECT Split_573_n1753_Split_574_n1754(net183_c1,net183);
INTERCONNECT Split_581_n1761_DFFT_187__FPB_n1367(net184_c1,net184);
INTERCONNECT Split_637_n1817_DFFT_193__FPB_n1373(net185_c1,net185);
INTERCONNECT Split_565_n1745_OR2T_48_n49(net186_c1,net186);
INTERCONNECT Split_557_n1737_AND2T_42_n43(net187_c1,net187);
INTERCONNECT Split_638_n1818_Split_640_n1820(net188_c1,net188);
INTERCONNECT Split_590_n1770_Split_591_n1771(net189_c1,net189);
INTERCONNECT Split_582_n1762_Split_583_n1763(net190_c1,net190);
INTERCONNECT Split_558_n1738_DFFT_243__FPB_n1423(net191_c1,net191);
INTERCONNECT Split_574_n1754_OR2T_98_n99(net192_c1,net192);
INTERCONNECT Split_566_n1746_DFFT_202__FPB_n1382(net193_c1,net193);
INTERCONNECT Split_591_n1771_OR2T_81_n82(net194_c1,net194);
INTERCONNECT Split_583_n1763_XOR2T_91_n92(net195_c1,net195);
INTERCONNECT Split_575_n1755_DFFT_400__FPB_n1580(net196_c1,net196);
INTERCONNECT Split_559_n1739_DFFT_150__FPB_n1330(net197_c1,net197);
INTERCONNECT Split_567_n1747_AND2T_66_n67(net198_c1,net198);
INTERCONNECT Split_639_n1819_OR2T_41_n42(net199_c1,net199);
INTERCONNECT Split_584_n1764_Split_586_n1766(net200_c1,net200);
INTERCONNECT Split_576_n1756_Split_578_n1758(net201_c1,net201);
INTERCONNECT Split_600_n1780_DFFT_383__FPB_n1563(net202_c1,net202);
INTERCONNECT Split_592_n1772_DFFT_434__FPB_n1614(net203_c1,net203);
INTERCONNECT Split_568_n1748_AND2T_88_n89(net204_c1,net204);
INTERCONNECT Split_593_n1773_Split_594_n1774(net205_c1,net205);
INTERCONNECT Split_577_n1757_DFFT_311__FPB_n1491(net206_c1,net206);
INTERCONNECT Split_601_n1781_AND2T_141_n142(net207_c1,net207);
INTERCONNECT Split_569_n1749_Split_570_n1750(net208_c1,net208);
INTERCONNECT Split_585_n1765_XOR2T_72_n73(net209_c1,net209);
INTERCONNECT Split_578_n1758_DFFT_482__FPB_n1662(net210_c1,net210);
INTERCONNECT Split_610_n1790_DFFT_207__FPB_n1387(net211_c1,net211);
INTERCONNECT Split_594_n1774_DFFT_264__FPB_n1444(net212_c1,net212);
INTERCONNECT Split_602_n1782_OR2T_111_n112(net213_c1,net213);
INTERCONNECT Split_586_n1766_DFFT_415__FPB_n1595(net214_c1,net214);
INTERCONNECT Split_611_n1791_Split_613_n1793(net215_c1,net215);
INTERCONNECT Split_579_n1759_Split_580_n1760(net216_c1,net216);
INTERCONNECT Split_603_n1783_XOR2T_128_n129(net217_c1,net217);
INTERCONNECT Split_587_n1767_DFFT_275__FPB_n1455(net218_c1,net218);
INTERCONNECT Split_595_n1775_DFFT_358__FPB_n1538(net219_c1,net219);
INTERCONNECT Split_588_n1768_DFFT_393__FPB_n1573(net220_c1,net220);
INTERCONNECT Split_604_n1784_XOR2T_128_n129(net221_c1,net221);
INTERCONNECT Split_596_n1776_AND2T_129_n130(net222_c1,net222);
INTERCONNECT Split_612_n1792_DFFT_148__FPB_n1328(net223_c1,net223);
INTERCONNECT Split_613_n1793_DFFT_167__FPB_n1347(net224_c1,net224);
INTERCONNECT Split_605_n1785_XOR2T_122_n123(net225_c1,net225);
INTERCONNECT Split_597_n1777_AND2T_118_n119(net226_c1,net226);
INTERCONNECT Split_589_n1769_DFFT_263__FPB_n1443(net227_c1,net227);
INTERCONNECT Split_614_n1794_Split_616_n1796(net228_c1,net228);
INTERCONNECT Split_606_n1786_AND2T_124_n125(net229_c1,net229);
INTERCONNECT Split_598_n1778_DFFT_386__FPB_n1566(net230_c1,net230);
INTERCONNECT Split_599_n1779_Split_600_n1780(net231_c1,net231);
INTERCONNECT Split_607_n1787_AND2T_132_n133(net232_c1,net232);
INTERCONNECT Split_615_n1795_OR2T_25_n25(net233_c1,net233);
INTERCONNECT Split_608_n1788_Split_610_n1790(net234_c1,net234);
INTERCONNECT Split_616_n1796_DFFT_156__FPB_n1336(net235_c1,net235);
INTERCONNECT Split_617_n1797_Split_619_n1799(net236_c1,net236);
INTERCONNECT Split_609_n1789_OR2T_30_n31(net237_c1,net237);
INTERCONNECT Split_618_n1798_AND2T_54_n55(net238_c1,net238);
INTERCONNECT Split_619_n1799_DFFT_282__FPB_n1462(net239_c1,net239);
INTERCONNECT Split_620_n1800_Split_621_n1801(net240_c1,net240);
INTERCONNECT Split_541_n1721_NOTT_139_n140(net241_c1,net241);
INTERCONNECT Split_621_n1801_AND2T_67_n68(net242_c1,net242);
INTERCONNECT Split_542_n1722_NOTT_58_n59(net243_c1,net243);
INTERCONNECT Split_550_n1730_NOTT_137_n138(net244_c1,net244);
INTERCONNECT Split_622_n1802_OR2T_73_n74(net245_c1,net245);
INTERCONNECT Split_630_n1810_OR2T_25_n25(net246_c1,net246);
INTERCONNECT Split_543_n1723_DFFT_229__FPB_n1409(net247_c1,net247);
INTERCONNECT Split_551_n1731_DFFT_254__FPB_n1434(net248_c1,net248);
INTERCONNECT Split_623_n1803_Split_624_n1804(net249_c1,net249);
INTERCONNECT Split_631_n1811_DFFT_153__FPB_n1333(net250_c1,net250);
INTERCONNECT Split_544_n1724_NOTT_56_n57(net251_c1,net251);
INTERCONNECT Split_552_n1732_DFFT_147__FPB_n148(net252_c1,net252);
INTERCONNECT Split_560_n1740_AND2T_28_n28(net253_c1,net253);
INTERCONNECT Split_624_n1804_OR2T_119_n120(net254_c1,net254);
INTERCONNECT Split_632_n1812_Split_633_n1813(net255_c1,net255);
INTERCONNECT Split_640_n1820_XOR2T_47_n48(net256_c1,net256);
INTERCONNECT Split_545_n1725_DFFT_252__FPB_n1432(net257_c1,net257);
INTERCONNECT Split_553_n1733_NOTT_138_n139(net258_c1,net258);
INTERCONNECT Split_561_n1741_OR2T_46_n47(net259_c1,net259);
INTERCONNECT Split_625_n1805_AND2T_131_n132(net260_c1,net260);
INTERCONNECT Split_633_n1813_NOTT_18_n18(net261_c1,net261);
INTERCONNECT Split_641_n1821_Split_642_n1822(net262_c1,net262);
INTERCONNECT Split_546_n1726_DFFT_186__FPB_n1366(net263_c1,net263);
INTERCONNECT Split_554_n1734_DFFT_299__FPB_n1479(net264_c1,net264);
INTERCONNECT Split_562_n1742_DFFT_477__FPB_n1657(net265_c1,net265);
INTERCONNECT Split_570_n1750_OR2T_45_n46(net266_c1,net266);
INTERCONNECT Split_626_n1806_Split_627_n1807(net267_c1,net267);
INTERCONNECT Split_634_n1814_DFFT_218__FPB_n1398(net268_c1,net268);
INTERCONNECT Split_642_n1822_XOR2T_62_n63(net269_c1,net269);
INTERCONNECT Split_547_n1727_NOTT_17_n17(net270_c1,net270);
INTERCONNECT Split_555_n1735_AND2T_19_n19(net271_c1,net271);
INTERCONNECT Split_563_n1743_AND2T_75_n76(net272_c1,net272);
INTERCONNECT Split_571_n1751_AND2T_140_n141(net273_c1,net273);
INTERCONNECT Split_627_n1807_OR2T_22_n22(net274_c1,net274);
INTERCONNECT Split_635_n1815_Split_636_n1816(net275_c1,net275);
INTERCONNECT Split_643_n1823_DFFT_190__FPB_n1370(net276_c1,net276);
INTERCONNECT Split_548_n1728_NOTT_136_n137(net277_c1,net277);
INTERCONNECT Split_556_n1736_DFFT_149__FPB_n1329(net278_c1,net278);
INTERCONNECT Split_564_n1744_OR2T_60_n61(net279_c1,net279);
INTERCONNECT Split_572_n1752_AND2T_53_n54(net280_c1,net280);
INTERCONNECT Split_580_n1760_AND2T_57_n58(net281_c1,net281);
INTERCONNECT Split_628_n1808_OR2T_30_n31(net282_c1,net282);
INTERCONNECT Split_636_n1816_NOTT_20_n20(net283_c1,net283);
INTERCONNECT Split_549_n1729_Split_550_n1730(net284_c1,net284);
INTERCONNECT Split_557_n1737_AND2T_27_n27(net285_c1,net285);
INTERCONNECT Split_565_n1745_OR2T_36_n37(net286_c1,net286);
INTERCONNECT Split_573_n1753_NOTT_107_n108(net287_c1,net287);
INTERCONNECT Split_581_n1761_XOR2T_62_n63(net288_c1,net288);
INTERCONNECT Split_629_n1809_Split_630_n1810(net289_c1,net289);
INTERCONNECT Split_637_n1817_OR2T_41_n42(net290_c1,net290);
INTERCONNECT Split_558_n1738_DFFT_179__FPB_n1359(net291_c1,net291);
INTERCONNECT Split_566_n1746_OR2T_37_n38(net292_c1,net292);
INTERCONNECT Split_574_n1754_AND2T_92_n93(net293_c1,net293);
INTERCONNECT Split_582_n1762_DFFT_277__FPB_n1457(net294_c1,net294);
INTERCONNECT Split_590_n1770_DFFT_344__FPB_n1524(net295_c1,net295);
INTERCONNECT Split_638_n1818_Split_639_n1819(net296_c1,net296);
INTERCONNECT Split_559_n1739_OR2T_40_n41(net297_c1,net297);
INTERCONNECT Split_567_n1747_AND2T_38_n39(net298_c1,net298);
INTERCONNECT Split_575_n1755_NOTT_55_n56(net299_c1,net299);
INTERCONNECT Split_583_n1763_AND2T_66_n67(net300_c1,net300);
INTERCONNECT Split_591_n1771_NOTT_77_n78(net301_c1,net301);
INTERCONNECT Split_639_n1819_NOTT_21_n21(net302_c1,net302);
INTERCONNECT Split_568_n1748_OR2T_52_n53(net303_c1,net303);
INTERCONNECT Split_576_n1756_Split_577_n1757(net304_c1,net304);
INTERCONNECT Split_584_n1764_Split_585_n1765(net305_c1,net305);
INTERCONNECT Split_592_n1772_OR2T_79_n80(net306_c1,net306);
INTERCONNECT Split_600_n1780_NOTT_101_n102(net307_c1,net307);
INTERCONNECT Split_569_n1749_OR2T_96_n97(net308_c1,net308);
INTERCONNECT Split_577_n1757_DFFT_286__FPB_n1466(net309_c1,net309);
INTERCONNECT Split_585_n1765_OR2T_71_n72(net310_c1,net310);
INTERCONNECT Split_593_n1773_DFFT_421__FPB_n1601(net311_c1,net311);
INTERCONNECT Split_601_n1781_AND2T_103_n104(net312_c1,net312);
INTERCONNECT Split_578_n1758_DFFT_369__FPB_n1549(net313_c1,net313);
INTERCONNECT Split_586_n1766_XOR2T_105_n106(net314_c1,net314);
INTERCONNECT Split_594_n1774_NOTT_110_n111(net315_c1,net315);
INTERCONNECT Split_602_n1782_OR2T_108_n109(net316_c1,net316);
INTERCONNECT Split_610_n1790_DFFT_168__FPB_n1348(net317_c1,net317);
INTERCONNECT Split_579_n1759_DFFT_335__FPB_n1515(net318_c1,net318);
INTERCONNECT Split_587_n1767_NOTT_104_n105(net319_c1,net319);
INTERCONNECT Split_595_n1775_NOTT_83_n84(net320_c1,net320);
INTERCONNECT Split_603_n1783_OR2T_113_n114(net321_c1,net321);
INTERCONNECT Split_611_n1791_Split_612_n1792(net322_c1,net322);
INTERCONNECT Split_588_n1768_DFFT_274__FPB_n1454(net323_c1,net323);
INTERCONNECT Split_596_n1776_OR2T_84_n85(net324_c1,net324);
INTERCONNECT Split_604_n1784_OR2T_113_n114(net325_c1,net325);
INTERCONNECT Split_612_n1792_OR2T_26_n26(net326_c1,net326);
INTERCONNECT Split_589_n1769_AND2T_78_n79(net327_c1,net327);
INTERCONNECT Split_597_n1777_AND2T_95_n96(net328_c1,net328);
INTERCONNECT Split_605_n1785_AND2T_114_n115(net329_c1,net329);
INTERCONNECT Split_613_n1793_DFFT_158__FPB_n1338(net330_c1,net330);
INTERCONNECT Split_598_n1778_AND2T_99_n100(net331_c1,net331);
INTERCONNECT Split_606_n1786_XOR2T_117_n118(net332_c1,net332);
INTERCONNECT Split_614_n1794_Split_615_n1795(net333_c1,net333);
INTERCONNECT Split_599_n1779_DFFT_397__FPB_n1577(net334_c1,net334);
INTERCONNECT Split_607_n1787_AND2T_126_n127(net335_c1,net335);
INTERCONNECT Split_615_n1795_OR2T_22_n22(net336_c1,net336);
INTERCONNECT Split_608_n1788_Split_609_n1789(net337_c1,net337);
INTERCONNECT Split_616_n1796_OR2T_39_n40(net338_c1,net338);
INTERCONNECT Split_609_n1789_AND2T_19_n19(net339_c1,net339);
INTERCONNECT Split_617_n1797_Split_618_n1798(net340_c1,net340);
INTERCONNECT Split_618_n1798_AND2T_33_n34(net341_c1,net341);
INTERCONNECT Split_619_n1799_DFFT_172__FPB_n1352(net342_c1,net342);
INTERCONNECT DFFT_220__FPB_n1400_DFFT_221__FPB_n1401(net343_c1,net343);
INTERCONNECT DFFT_221__FPB_n1401_DFFT_222__FPB_n1402(net344_c1,net344);
INTERCONNECT DFFT_230__FPB_n1410_DFFT_231__FPB_n1411(net345_c1,net345);
INTERCONNECT DFFT_222__FPB_n1402_DFFT_223__FPB_n1403(net346_c1,net346);
INTERCONNECT DFFT_150__FPB_n1330_Split_HOLD_1685(net347_c1,net347);
INTERCONNECT DFFT_231__FPB_n1411_DFFT_232__FPB_n1412(net348_c1,net348);
INTERCONNECT DFFT_223__FPB_n1403_DFFT_224__FPB_n1404(net349_c1,net349);
INTERCONNECT DFFT_151__FPB_n1331_AND2T_29_n30(net350_c1,net350);
INTERCONNECT DFFT_320__FPB_n1500_DFFT_321__FPB_n1501(net351_c1,net351);
INTERCONNECT DFFT_240__FPB_n1420_DFFT_241__FPB_n1421(net352_c1,net352);
INTERCONNECT DFFT_232__FPB_n1412_Split_HOLD_1678(net353_c1,net353);
INTERCONNECT DFFT_224__FPB_n1404_DFFT_225__FPB_n1405(net354_c1,net354);
INTERCONNECT DFFT_160__FPB_n1340_DFFT_161__FPB_n1341(net355_c1,net355);
INTERCONNECT DFFT_152__FPB_n1332_OR2T_31_n32(net356_c1,net356);
INTERCONNECT DFFT_321__FPB_n1501_DFFT_322__FPB_n1502(net357_c1,net357);
INTERCONNECT DFFT_241__FPB_n1421_DFFT_242__FPB_n1422(net358_c1,net358);
INTERCONNECT DFFT_233__FPB_n1413_DFFT_234__FPB_n1414(net359_c1,net359);
INTERCONNECT DFFT_225__FPB_n1405_DFFT_226__FPB_n1406(net360_c1,net360);
INTERCONNECT DFFT_153__FPB_n1333_DFFT_154__FPB_n1334(net361_c1,net361);
INTERCONNECT DFFT_161__FPB_n1341_OR2T_37_n38(net362_c1,net362);
INTERCONNECT DFFT_330__FPB_n1510_Split_HOLD_1676(net363_c1,net363);
INTERCONNECT DFFT_322__FPB_n1502_DFFT_323__FPB_n1503(net364_c1,net364);
INTERCONNECT DFFT_250__FPB_n1430_DFFT_251__FPB_n1431(net365_c1,net365);
INTERCONNECT DFFT_234__FPB_n1414_DFFT_235__FPB_n1415(net366_c1,net366);
INTERCONNECT DFFT_226__FPB_n1406_DFFT_227__FPB_n1407(net367_c1,net367);
INTERCONNECT DFFT_170__FPB_n1350_DFFT_171__FPB_n1351(net368_c1,net368);
INTERCONNECT DFFT_162__FPB_n1342_DFFT_163__FPB_n1343(net369_c1,net369);
INTERCONNECT DFFT_154__FPB_n1334_DFFT_155__FPB_n1335(net370_c1,net370);
INTERCONNECT DFFT_242__FPB_n1422_AND2T_76_n77(net371_c1,net371);
INTERCONNECT DFFT_331__FPB_n1511_DFFT_332__FPB_n1512(net372_c1,net372);
INTERCONNECT DFFT_323__FPB_n1503_DFFT_324__FPB_n1504(net373_c1,net373);
INTERCONNECT DFFT_243__FPB_n1423_DFFT_244__FPB_n1424(net374_c1,net374);
INTERCONNECT DFFT_235__FPB_n1415_DFFT_236__FPB_n1416(net375_c1,net375);
INTERCONNECT DFFT_227__FPB_n1407_DFFT_228__FPB_n1408(net376_c1,net376);
INTERCONNECT DFFT_163__FPB_n1343_DFFT_164__FPB_n1344(net377_c1,net377);
INTERCONNECT DFFT_251__FPB_n1431_OR2T_79_n80(net378_c1,net378);
INTERCONNECT DFFT_171__FPB_n1351_XOR2T_44_n45(net379_c1,net379);
INTERCONNECT DFFT_155__FPB_n1335_AND2T_35_n36(net380_c1,net380);
INTERCONNECT DFFT_340__FPB_n1520_DFFT_341__FPB_n1521(net381_c1,net381);
INTERCONNECT DFFT_332__FPB_n1512_DFFT_333__FPB_n1513(net382_c1,net382);
INTERCONNECT DFFT_260__FPB_n1440_DFFT_261__FPB_n1441(net383_c1,net383);
INTERCONNECT DFFT_252__FPB_n1432_DFFT_253__FPB_n1433(net384_c1,net384);
INTERCONNECT DFFT_244__FPB_n1424_DFFT_245__FPB_n1425(net385_c1,net385);
INTERCONNECT DFFT_236__FPB_n1416_DFFT_237__FPB_n1417(net386_c1,net386);
INTERCONNECT DFFT_172__FPB_n1352_DFFT_173__FPB_n1353(net387_c1,net387);
INTERCONNECT DFFT_164__FPB_n1344_DFFT_165__FPB_n1345(net388_c1,net388);
INTERCONNECT DFFT_156__FPB_n1336_DFFT_157__FPB_n1337(net389_c1,net389);
INTERCONNECT DFFT_420__FPB_n1600_AND2T_126_n127(net390_c1,net390);
INTERCONNECT DFFT_324__FPB_n1504_AND2T_103_n104(net391_c1,net391);
INTERCONNECT DFFT_228__FPB_n1408_XOR2T_72_n73(net392_c1,net392);
INTERCONNECT DFFT_180__FPB_n1360_AND2T_49_n50(net393_c1,net393);
INTERCONNECT DFFT_148__FPB_n1328_AND2T_23_n23(net394_c1,net394);
INTERCONNECT DFFT_421__FPB_n1601_DFFT_422__FPB_n1602(net395_c1,net395);
INTERCONNECT DFFT_341__FPB_n1521_DFFT_342__FPB_n1522(net396_c1,net396);
INTERCONNECT DFFT_333__FPB_n1513_DFFT_334__FPB_n1514(net397_c1,net397);
INTERCONNECT DFFT_325__FPB_n1505_DFFT_326__FPB_n1506(net398_c1,net398);
INTERCONNECT DFFT_261__FPB_n1441_DFFT_262__FPB_n1442(net399_c1,net399);
INTERCONNECT DFFT_245__FPB_n1425_DFFT_246__FPB_n1426(net400_c1,net400);
INTERCONNECT DFFT_229__FPB_n1409_DFFT_230__FPB_n1410(net401_c1,net401);
INTERCONNECT DFFT_181__FPB_n1361_DFFT_182__FPB_n1362(net402_c1,net402);
INTERCONNECT DFFT_173__FPB_n1353_DFFT_174__FPB_n1354(net403_c1,net403);
INTERCONNECT DFFT_253__FPB_n1433_OR2T_80_n81(net404_c1,net404);
INTERCONNECT DFFT_237__FPB_n1417_OR2T_73_n74(net405_c1,net405);
INTERCONNECT DFFT_165__FPB_n1345_AND2T_38_n39(net406_c1,net406);
INTERCONNECT DFFT_157__FPB_n1337_OR2T_36_n37(net407_c1,net407);
INTERCONNECT DFFT_149__FPB_n1329_AND2T_24_n24(net408_c1,net408);
INTERCONNECT DFFT_422__FPB_n1602_DFFT_423__FPB_n1603(net409_c1,net409);
INTERCONNECT DFFT_350__FPB_n1530_DFFT_351__FPB_n1531(net410_c1,net410);
INTERCONNECT DFFT_342__FPB_n1522_Split_HOLD_1673(net411_c1,net411);
INTERCONNECT DFFT_326__FPB_n1506_DFFT_327__FPB_n1507(net412_c1,net412);
INTERCONNECT DFFT_270__FPB_n1450_DFFT_271__FPB_n1451(net413_c1,net413);
INTERCONNECT DFFT_254__FPB_n1434_DFFT_255__FPB_n1435(net414_c1,net414);
INTERCONNECT DFFT_246__FPB_n1426_DFFT_247__FPB_n1427(net415_c1,net415);
INTERCONNECT DFFT_190__FPB_n1370_DFFT_191__FPB_n1371(net416_c1,net416);
INTERCONNECT DFFT_182__FPB_n1362_DFFT_183__FPB_n1363(net417_c1,net417);
INTERCONNECT DFFT_158__FPB_n1338_DFFT_159__FPB_n1339(net418_c1,net418);
INTERCONNECT DFFT_430__FPB_n1610_OR2T_130_n131(net419_c1,net419);
INTERCONNECT DFFT_334__FPB_n1514_XOR2T_105_n106(net420_c1,net420);
INTERCONNECT DFFT_262__FPB_n1442_OR2T_81_n82(net421_c1,net421);
INTERCONNECT DFFT_238__FPB_n1418_AND2T_75_n76(net422_c1,net422);
INTERCONNECT DFFT_174__FPB_n1354_OR2T_45_n46(net423_c1,net423);
INTERCONNECT DFFT_166__FPB_n1346_OR2T_39_n40(net424_c1,net424);
INTERCONNECT DFFT_431__FPB_n1611_DFFT_432__FPB_n1612(net425_c1,net425);
INTERCONNECT DFFT_423__FPB_n1603_DFFT_424__FPB_n1604(net426_c1,net426);
INTERCONNECT DFFT_351__FPB_n1531_DFFT_352__FPB_n1532(net427_c1,net427);
INTERCONNECT DFFT_335__FPB_n1515_DFFT_336__FPB_n1516(net428_c1,net428);
INTERCONNECT DFFT_327__FPB_n1507_DFFT_328__FPB_n1508(net429_c1,net429);
INTERCONNECT DFFT_271__FPB_n1451_DFFT_272__FPB_n1452(net430_c1,net430);
INTERCONNECT DFFT_255__FPB_n1435_DFFT_256__FPB_n1436(net431_c1,net431);
INTERCONNECT DFFT_247__FPB_n1427_DFFT_248__FPB_n1428(net432_c1,net432);
INTERCONNECT DFFT_239__FPB_n1419_DFFT_240__FPB_n1420(net433_c1,net433);
INTERCONNECT DFFT_183__FPB_n1363_DFFT_184__FPB_n1364(net434_c1,net434);
INTERCONNECT DFFT_175__FPB_n1355_DFFT_176__FPB_n1356(net435_c1,net435);
INTERCONNECT DFFT_159__FPB_n1339_DFFT_160__FPB_n1340(net436_c1,net436);
INTERCONNECT DFFT_343__FPB_n1523_AND2T_106_n107(net437_c1,net437);
INTERCONNECT DFFT_263__FPB_n1443_AND2T_82_n83(net438_c1,net438);
INTERCONNECT DFFT_191__FPB_n1371_OR2T_60_n61(net439_c1,net439);
INTERCONNECT DFFT_167__FPB_n1347_OR2T_40_n41(net440_c1,net440);
INTERCONNECT DFFT_520__FPB_n1700_DFFT_521__FPB_n1701(net441_c1,net441);
INTERCONNECT DFFT_432__FPB_n1612_DFFT_433__FPB_n1613(net442_c1,net442);
INTERCONNECT DFFT_424__FPB_n1604_DFFT_425__FPB_n1605(net443_c1,net443);
INTERCONNECT DFFT_360__FPB_n1540_DFFT_361__FPB_n1541(net444_c1,net444);
INTERCONNECT DFFT_352__FPB_n1532_DFFT_353__FPB_n1533(net445_c1,net445);
INTERCONNECT DFFT_344__FPB_n1524_DFFT_345__FPB_n1525(net446_c1,net446);
INTERCONNECT DFFT_336__FPB_n1516_DFFT_337__FPB_n1517(net447_c1,net447);
INTERCONNECT DFFT_328__FPB_n1508_DFFT_329__FPB_n1509(net448_c1,net448);
INTERCONNECT DFFT_280__FPB_n1460_DFFT_281__FPB_n1461(net449_c1,net449);
INTERCONNECT DFFT_264__FPB_n1444_DFFT_265__FPB_n1445(net450_c1,net450);
INTERCONNECT DFFT_256__FPB_n1436_DFFT_257__FPB_n1437(net451_c1,net451);
INTERCONNECT DFFT_248__FPB_n1428_DFFT_249__FPB_n1429(net452_c1,net452);
INTERCONNECT DFFT_184__FPB_n1364_DFFT_185__FPB_n1365(net453_c1,net453);
INTERCONNECT DFFT_176__FPB_n1356_Split_HOLD_1672(net454_c1,net454);
INTERCONNECT DFFT_168__FPB_n1348_DFFT_169__FPB_n1349(net455_c1,net455);
INTERCONNECT DFFT_440__FPB_n1620_AND2T_132_n133(net456_c1,net456);
INTERCONNECT DFFT_272__FPB_n1452_OR2T_84_n85(net457_c1,net457);
INTERCONNECT DFFT_200__FPB_n1380_XOR2T_65_n66(net458_c1,net458);
INTERCONNECT DFFT_192__FPB_n1372_AND2T_61_n62(net459_c1,net459);
INTERCONNECT DFFT_521__FPB_n1701_DFFT_522__FPB_n1702(net460_c1,net460);
INTERCONNECT DFFT_441__FPB_n1621_DFFT_442__FPB_n1622(net461_c1,net461);
INTERCONNECT DFFT_425__FPB_n1605_DFFT_426__FPB_n1606(net462_c1,net462);
INTERCONNECT DFFT_361__FPB_n1541_DFFT_362__FPB_n1542(net463_c1,net463);
INTERCONNECT DFFT_353__FPB_n1533_DFFT_354__FPB_n1534(net464_c1,net464);
INTERCONNECT DFFT_337__FPB_n1517_DFFT_338__FPB_n1518(net465_c1,net465);
INTERCONNECT DFFT_329__FPB_n1509_DFFT_330__FPB_n1510(net466_c1,net466);
INTERCONNECT DFFT_265__FPB_n1445_DFFT_266__FPB_n1446(net467_c1,net467);
INTERCONNECT DFFT_257__FPB_n1437_DFFT_258__FPB_n1438(net468_c1,net468);
INTERCONNECT DFFT_249__FPB_n1429_DFFT_250__FPB_n1430(net469_c1,net469);
INTERCONNECT DFFT_193__FPB_n1373_DFFT_194__FPB_n1374(net470_c1,net470);
INTERCONNECT DFFT_169__FPB_n1349_DFFT_170__FPB_n1350(net471_c1,net471);
INTERCONNECT DFFT_433__FPB_n1613_AND2T_131_n132(net472_c1,net472);
INTERCONNECT DFFT_345__FPB_n1525_OR2T_108_n109(net473_c1,net473);
INTERCONNECT DFFT_281__FPB_n1461_XOR2T_89_n90(net474_c1,net474);
INTERCONNECT DFFT_273__FPB_n1453_AND2T_85_n86(net475_c1,net475);
INTERCONNECT DFFT_201__FPB_n1381_AND2T_67_n68(net476_c1,net476);
INTERCONNECT DFFT_185__FPB_n1365_AND2T_53_n54(net477_c1,net477);
INTERCONNECT DFFT_177__FPB_n1357_OR2T_46_n47(net478_c1,net478);
INTERCONNECT DFFT_530__FPB_n1710_DFFT_531__FPB_n1711(net479_c1,net479);
INTERCONNECT DFFT_522__FPB_n1702_DFFT_523__FPB_n1703(net480_c1,net480);
INTERCONNECT DFFT_450__FPB_n1630_DFFT_451__FPB_n1631(net481_c1,net481);
INTERCONNECT DFFT_442__FPB_n1622_DFFT_443__FPB_n1623(net482_c1,net482);
INTERCONNECT DFFT_434__FPB_n1614_DFFT_435__FPB_n1615(net483_c1,net483);
INTERCONNECT DFFT_426__FPB_n1606_Split_HOLD_1670(net484_c1,net484);
INTERCONNECT DFFT_370__FPB_n1550_DFFT_371__FPB_n1551(net485_c1,net485);
INTERCONNECT DFFT_362__FPB_n1542_DFFT_363__FPB_n1543(net486_c1,net486);
INTERCONNECT DFFT_354__FPB_n1534_DFFT_355__FPB_n1535(net487_c1,net487);
INTERCONNECT DFFT_346__FPB_n1526_DFFT_347__FPB_n1527(net488_c1,net488);
INTERCONNECT DFFT_338__FPB_n1518_DFFT_339__FPB_n1519(net489_c1,net489);
INTERCONNECT DFFT_290__FPB_n1470_Split_HOLD_1669(net490_c1,net490);
INTERCONNECT DFFT_282__FPB_n1462_DFFT_283__FPB_n1463(net491_c1,net491);
INTERCONNECT DFFT_266__FPB_n1446_DFFT_267__FPB_n1447(net492_c1,net492);
INTERCONNECT DFFT_258__FPB_n1438_DFFT_259__FPB_n1439(net493_c1,net493);
INTERCONNECT DFFT_210__FPB_n1390_DFFT_211__FPB_n1391(net494_c1,net494);
INTERCONNECT DFFT_202__FPB_n1382_DFFT_203__FPB_n1383(net495_c1,net495);
INTERCONNECT DFFT_194__FPB_n1374_Split_HOLD_1668(net496_c1,net496);
INTERCONNECT DFFT_274__FPB_n1454_OR2T_86_n87(net497_c1,net497);
INTERCONNECT DFFT_186__FPB_n1366_AND2T_54_n55(net498_c1,net498);
INTERCONNECT DFFT_178__FPB_n1358_OR2T_48_n49(net499_c1,net499);
INTERCONNECT DFFT_531__FPB_n1711_DFFT_532__FPB_n1712(net500_c1,net500);
INTERCONNECT DFFT_523__FPB_n1703_DFFT_524__FPB_n1704(net501_c1,net501);
INTERCONNECT DFFT_451__FPB_n1631_DFFT_452__FPB_n1632(net502_c1,net502);
INTERCONNECT DFFT_443__FPB_n1623_DFFT_444__FPB_n1624(net503_c1,net503);
INTERCONNECT DFFT_435__FPB_n1615_DFFT_436__FPB_n1616(net504_c1,net504);
INTERCONNECT DFFT_427__FPB_n1607_DFFT_428__FPB_n1608(net505_c1,net505);
INTERCONNECT DFFT_371__FPB_n1551_DFFT_372__FPB_n1552(net506_c1,net506);
INTERCONNECT DFFT_363__FPB_n1543_DFFT_364__FPB_n1544(net507_c1,net507);
INTERCONNECT DFFT_355__FPB_n1535_DFFT_356__FPB_n1536(net508_c1,net508);
INTERCONNECT DFFT_347__FPB_n1527_DFFT_348__FPB_n1528(net509_c1,net509);
INTERCONNECT DFFT_339__FPB_n1519_DFFT_340__FPB_n1520(net510_c1,net510);
INTERCONNECT DFFT_291__FPB_n1471_DFFT_292__FPB_n1472(net511_c1,net511);
INTERCONNECT DFFT_283__FPB_n1463_DFFT_284__FPB_n1464(net512_c1,net512);
INTERCONNECT DFFT_275__FPB_n1455_DFFT_276__FPB_n1456(net513_c1,net513);
INTERCONNECT DFFT_267__FPB_n1447_DFFT_268__FPB_n1448(net514_c1,net514);
INTERCONNECT DFFT_259__FPB_n1439_DFFT_260__FPB_n1440(net515_c1,net515);
INTERCONNECT DFFT_211__FPB_n1391_DFFT_212__FPB_n1392(net516_c1,net516);
INTERCONNECT DFFT_203__FPB_n1383_DFFT_204__FPB_n1384(net517_c1,net517);
INTERCONNECT DFFT_187__FPB_n1367_DFFT_188__FPB_n1368(net518_c1,net518);
INTERCONNECT DFFT_179__FPB_n1359_DFFT_180__FPB_n1360(net519_c1,net519);
INTERCONNECT DFFT_195__FPB_n1375_OR2T_63_n64(net520_c1,net520);
INTERCONNECT DFFT_532__FPB_n1712_DFFT_533__FPB_n1713(net521_c1,net521);
INTERCONNECT DFFT_524__FPB_n1704_DFFT_525__FPB_n1705(net522_c1,net522);
INTERCONNECT DFFT_460__FPB_n1640_DFFT_461__FPB_n1641(net523_c1,net523);
INTERCONNECT DFFT_452__FPB_n1632_DFFT_453__FPB_n1633(net524_c1,net524);
INTERCONNECT DFFT_444__FPB_n1624_DFFT_445__FPB_n1625(net525_c1,net525);
INTERCONNECT DFFT_436__FPB_n1616_DFFT_437__FPB_n1617(net526_c1,net526);
INTERCONNECT DFFT_428__FPB_n1608_DFFT_429__FPB_n1609(net527_c1,net527);
INTERCONNECT DFFT_380__FPB_n1560_DFFT_381__FPB_n1561(net528_c1,net528);
INTERCONNECT DFFT_372__FPB_n1552_DFFT_373__FPB_n1553(net529_c1,net529);
INTERCONNECT DFFT_364__FPB_n1544_DFFT_365__FPB_n1545(net530_c1,net530);
INTERCONNECT DFFT_356__FPB_n1536_DFFT_357__FPB_n1537(net531_c1,net531);
INTERCONNECT DFFT_348__FPB_n1528_DFFT_349__FPB_n1529(net532_c1,net532);
INTERCONNECT DFFT_300__FPB_n1480_DFFT_301__FPB_n1481(net533_c1,net533);
INTERCONNECT DFFT_292__FPB_n1472_DFFT_293__FPB_n1473(net534_c1,net534);
INTERCONNECT DFFT_268__FPB_n1448_DFFT_269__FPB_n1449(net535_c1,net535);
INTERCONNECT DFFT_212__FPB_n1392_DFFT_213__FPB_n1393(net536_c1,net536);
INTERCONNECT DFFT_204__FPB_n1384_DFFT_205__FPB_n1385(net537_c1,net537);
INTERCONNECT DFFT_196__FPB_n1376_DFFT_197__FPB_n1377(net538_c1,net538);
INTERCONNECT DFFT_188__FPB_n1368_DFFT_189__FPB_n1369(net539_c1,net539);
INTERCONNECT DFFT_284__FPB_n1464_OR2T_90_n91(net540_c1,net540);
INTERCONNECT DFFT_276__FPB_n1456_AND2T_87_n88(net541_c1,net541);
INTERCONNECT DFFT_533__FPB_n1713_DFFT_534__FPB_n1714(net542_c1,net542);
INTERCONNECT DFFT_525__FPB_n1705_DFFT_526__FPB_n1706(net543_c1,net543);
INTERCONNECT DFFT_461__FPB_n1641_DFFT_462__FPB_n1642(net544_c1,net544);
INTERCONNECT DFFT_453__FPB_n1633_DFFT_454__FPB_n1634(net545_c1,net545);
INTERCONNECT DFFT_445__FPB_n1625_DFFT_446__FPB_n1626(net546_c1,net546);
INTERCONNECT DFFT_437__FPB_n1617_DFFT_438__FPB_n1618(net547_c1,net547);
INTERCONNECT DFFT_381__FPB_n1561_DFFT_382__FPB_n1562(net548_c1,net548);
INTERCONNECT DFFT_373__FPB_n1553_DFFT_374__FPB_n1554(net549_c1,net549);
INTERCONNECT DFFT_365__FPB_n1545_DFFT_366__FPB_n1546(net550_c1,net550);
INTERCONNECT DFFT_349__FPB_n1529_DFFT_350__FPB_n1530(net551_c1,net551);
INTERCONNECT DFFT_301__FPB_n1481_DFFT_302__FPB_n1482(net552_c1,net552);
INTERCONNECT DFFT_269__FPB_n1449_Split_HOLD_1667(net553_c1,net553);
INTERCONNECT DFFT_213__FPB_n1393_DFFT_214__FPB_n1394(net554_c1,net554);
INTERCONNECT DFFT_197__FPB_n1377_DFFT_198__FPB_n1378(net555_c1,net555);
INTERCONNECT DFFT_429__FPB_n1609_AND2T_129_n130(net556_c1,net556);
INTERCONNECT DFFT_357__FPB_n1537_AND2T_109_n110(net557_c1,net557);
INTERCONNECT DFFT_293__FPB_n1473_AND2T_95_n96(net558_c1,net558);
INTERCONNECT DFFT_285__FPB_n1465_XOR2T_93_n94(net559_c1,net559);
INTERCONNECT DFFT_277__FPB_n1457_AND2T_88_n89(net560_c1,net560);
INTERCONNECT DFFT_205__FPB_n1385_OR2T_68_n69(net561_c1,net561);
INTERCONNECT DFFT_189__FPB_n1369_AND2T_59_n60(net562_c1,net562);
INTERCONNECT DFFT_534__FPB_n1714_DFFT_535__FPB_n1715(net563_c1,net563);
INTERCONNECT DFFT_526__FPB_n1706_DFFT_527_Q2(net564_c1,net564);
INTERCONNECT DFFT_470__FPB_n1650_DFFT_471__FPB_n1651(net565_c1,net565);
INTERCONNECT DFFT_462__FPB_n1642_DFFT_463__FPB_n1643(net566_c1,net566);
INTERCONNECT DFFT_454__FPB_n1634_DFFT_455__FPB_n1635(net567_c1,net567);
INTERCONNECT DFFT_446__FPB_n1626_DFFT_447__FPB_n1627(net568_c1,net568);
INTERCONNECT DFFT_438__FPB_n1618_DFFT_439__FPB_n1619(net569_c1,net569);
INTERCONNECT DFFT_390__FPB_n1570_DFFT_391__FPB_n1571(net570_c1,net570);
INTERCONNECT DFFT_374__FPB_n1554_DFFT_375__FPB_n1555(net571_c1,net571);
INTERCONNECT DFFT_302__FPB_n1482_DFFT_303__FPB_n1483(net572_c1,net572);
INTERCONNECT DFFT_294__FPB_n1474_DFFT_295__FPB_n1475(net573_c1,net573);
INTERCONNECT DFFT_286__FPB_n1466_DFFT_287__FPB_n1467(net574_c1,net574);
INTERCONNECT DFFT_278__FPB_n1458_DFFT_279__FPB_n1459(net575_c1,net575);
INTERCONNECT DFFT_214__FPB_n1394_DFFT_215__FPB_n1395(net576_c1,net576);
INTERCONNECT DFFT_198__FPB_n1378_DFFT_199__FPB_n1379(net577_c1,net577);
INTERCONNECT DFFT_382__FPB_n1562_AND2T_116_n117(net578_c1,net578);
INTERCONNECT DFFT_366__FPB_n1546_AND2T_112_n113(net579_c1,net579);
INTERCONNECT DFFT_358__FPB_n1538_OR2T_111_n112(net580_c1,net580);
INTERCONNECT DFFT_310__FPB_n1490_OR2T_102_n103(net581_c1,net581);
INTERCONNECT DFFT_206__FPB_n1386_AND2T_69_n70(net582_c1,net582);
INTERCONNECT DFFT_535__FPB_n1715_DFFT_536__FPB_n1716(net583_c1,net583);
INTERCONNECT DFFT_471__FPB_n1651_DFFT_472__FPB_n1652(net584_c1,net584);
INTERCONNECT DFFT_463__FPB_n1643_DFFT_464__FPB_n1644(net585_c1,net585);
INTERCONNECT DFFT_455__FPB_n1635_DFFT_456__FPB_n1636(net586_c1,net586);
INTERCONNECT DFFT_447__FPB_n1627_DFFT_448__FPB_n1628(net587_c1,net587);
INTERCONNECT DFFT_439__FPB_n1619_DFFT_440__FPB_n1620(net588_c1,net588);
INTERCONNECT DFFT_391__FPB_n1571_DFFT_392__FPB_n1572(net589_c1,net589);
INTERCONNECT DFFT_383__FPB_n1563_DFFT_384__FPB_n1564(net590_c1,net590);
INTERCONNECT DFFT_375__FPB_n1555_DFFT_376__FPB_n1556(net591_c1,net591);
INTERCONNECT DFFT_359__FPB_n1539_DFFT_360__FPB_n1540(net592_c1,net592);
INTERCONNECT DFFT_311__FPB_n1491_DFFT_312__FPB_n1492(net593_c1,net593);
INTERCONNECT DFFT_303__FPB_n1483_DFFT_304__FPB_n1484(net594_c1,net594);
INTERCONNECT DFFT_287__FPB_n1467_DFFT_288__FPB_n1468(net595_c1,net595);
INTERCONNECT DFFT_279__FPB_n1459_DFFT_280__FPB_n1460(net596_c1,net596);
INTERCONNECT DFFT_215__FPB_n1395_Split_HOLD_1679(net597_c1,net597);
INTERCONNECT DFFT_207__FPB_n1387_DFFT_208__FPB_n1388(net598_c1,net598);
INTERCONNECT DFFT_199__FPB_n1379_DFFT_200__FPB_n1380(net599_c1,net599);
INTERCONNECT DFFT_367__FPB_n1547_AND2T_114_n115(net600_c1,net600);
INTERCONNECT DFFT_295__FPB_n1475_OR2T_96_n97(net601_c1,net601);
INTERCONNECT DFFT_536__FPB_n1716_DFFT_537__FPB_n1717(net602_c1,net602);
INTERCONNECT DFFT_528__FPB_n1708_DFFT_529__FPB_n1709(net603_c1,net603);
INTERCONNECT DFFT_480__FPB_n1660_DFFT_481__FPB_n1661(net604_c1,net604);
INTERCONNECT DFFT_472__FPB_n1652_DFFT_473__FPB_n1653(net605_c1,net605);
INTERCONNECT DFFT_464__FPB_n1644_DFFT_465__FPB_n1645(net606_c1,net606);
INTERCONNECT DFFT_456__FPB_n1636_Split_HOLD_1684(net607_c1,net607);
INTERCONNECT DFFT_448__FPB_n1628_DFFT_449__FPB_n1629(net608_c1,net608);
INTERCONNECT DFFT_400__FPB_n1580_DFFT_401__FPB_n1581(net609_c1,net609);
INTERCONNECT DFFT_384__FPB_n1564_Split_HOLD_1683(net610_c1,net610);
INTERCONNECT DFFT_376__FPB_n1556_DFFT_377__FPB_n1557(net611_c1,net611);
INTERCONNECT DFFT_312__FPB_n1492_DFFT_313__FPB_n1493(net612_c1,net612);
INTERCONNECT DFFT_304__FPB_n1484_DFFT_305__FPB_n1485(net613_c1,net613);
INTERCONNECT DFFT_296__FPB_n1476_DFFT_297__FPB_n1477(net614_c1,net614);
INTERCONNECT DFFT_288__FPB_n1468_DFFT_289__FPB_n1469(net615_c1,net615);
INTERCONNECT DFFT_216__FPB_n1396_DFFT_217__FPB_n1397(net616_c1,net616);
INTERCONNECT DFFT_208__FPB_n1388_DFFT_209__FPB_n1389(net617_c1,net617);
INTERCONNECT DFFT_392__FPB_n1572_OR2T_119_n120(net618_c1,net618);
INTERCONNECT DFFT_368__FPB_n1548_OR2T_115_n116(net619_c1,net619);
INTERCONNECT DFFT_537__FPB_n1717_DFFT_538_Q1(net620_c1,net620);
INTERCONNECT DFFT_529__FPB_n1709_DFFT_530__FPB_n1710(net621_c1,net621);
INTERCONNECT DFFT_473__FPB_n1653_DFFT_474__FPB_n1654(net622_c1,net622);
INTERCONNECT DFFT_465__FPB_n1645_DFFT_466__FPB_n1646(net623_c1,net623);
INTERCONNECT DFFT_457__FPB_n1637_DFFT_458__FPB_n1638(net624_c1,net624);
INTERCONNECT DFFT_449__FPB_n1629_DFFT_450__FPB_n1630(net625_c1,net625);
INTERCONNECT DFFT_401__FPB_n1581_DFFT_402__FPB_n1582(net626_c1,net626);
INTERCONNECT DFFT_377__FPB_n1557_DFFT_378__FPB_n1558(net627_c1,net627);
INTERCONNECT DFFT_369__FPB_n1549_DFFT_370__FPB_n1550(net628_c1,net628);
INTERCONNECT DFFT_313__FPB_n1493_DFFT_314__FPB_n1494(net629_c1,net629);
INTERCONNECT DFFT_305__FPB_n1485_DFFT_306__FPB_n1486(net630_c1,net630);
INTERCONNECT DFFT_297__FPB_n1477_Split_HOLD_1682(net631_c1,net631);
INTERCONNECT DFFT_289__FPB_n1469_DFFT_290__FPB_n1470(net632_c1,net632);
INTERCONNECT DFFT_209__FPB_n1389_Split_HOLD_1677(net633_c1,net633);
INTERCONNECT DFFT_481__FPB_n1661_AND2T_140_n141(net634_c1,net634);
INTERCONNECT DFFT_393__FPB_n1573_XOR2T_122_n123(net635_c1,net635);
INTERCONNECT DFFT_385__FPB_n1565_XOR2T_117_n118(net636_c1,net636);
INTERCONNECT DFFT_217__FPB_n1397_OR2T_71_n72(net637_c1,net637);
INTERCONNECT DFFT_490__FPB_n1670_DFFT_491__FPB_n1671(net638_c1,net638);
INTERCONNECT DFFT_482__FPB_n1662_DFFT_483__FPB_n1663(net639_c1,net639);
INTERCONNECT DFFT_474__FPB_n1654_DFFT_475__FPB_n1655(net640_c1,net640);
INTERCONNECT DFFT_466__FPB_n1646_DFFT_467__FPB_n1647(net641_c1,net641);
INTERCONNECT DFFT_458__FPB_n1638_DFFT_459__FPB_n1639(net642_c1,net642);
INTERCONNECT DFFT_410__FPB_n1590_DFFT_411__FPB_n1591(net643_c1,net643);
INTERCONNECT DFFT_402__FPB_n1582_DFFT_403__FPB_n1583(net644_c1,net644);
INTERCONNECT DFFT_394__FPB_n1574_DFFT_395__FPB_n1575(net645_c1,net645);
INTERCONNECT DFFT_378__FPB_n1558_DFFT_379__FPB_n1559(net646_c1,net646);
INTERCONNECT DFFT_314__FPB_n1494_DFFT_315__FPB_n1495(net647_c1,net647);
INTERCONNECT DFFT_306__FPB_n1486_DFFT_307__FPB_n1487(net648_c1,net648);
INTERCONNECT DFFT_218__FPB_n1398_DFFT_219__FPB_n1399(net649_c1,net649);
INTERCONNECT DFFT_386__FPB_n1566_AND2T_118_n119(net650_c1,net650);
INTERCONNECT DFFT_298__FPB_n1478_OR2T_98_n99(net651_c1,net651);
INTERCONNECT DFFT_539__FPB_n1719_DFFT_540_Q0(net652_c1,net652);
INTERCONNECT DFFT_491__FPB_n1671_DFFT_492__FPB_n1672(net653_c1,net653);
INTERCONNECT DFFT_483__FPB_n1663_DFFT_484__FPB_n1664(net654_c1,net654);
INTERCONNECT DFFT_475__FPB_n1655_DFFT_476__FPB_n1656(net655_c1,net655);
INTERCONNECT DFFT_467__FPB_n1647_DFFT_468__FPB_n1648(net656_c1,net656);
INTERCONNECT DFFT_411__FPB_n1591_DFFT_412__FPB_n1592(net657_c1,net657);
INTERCONNECT DFFT_403__FPB_n1583_Split_HOLD_1675(net658_c1,net658);
INTERCONNECT DFFT_395__FPB_n1575_DFFT_396__FPB_n1576(net659_c1,net659);
INTERCONNECT DFFT_387__FPB_n1567_Split_HOLD_1681(net660_c1,net660);
INTERCONNECT DFFT_379__FPB_n1559_DFFT_380__FPB_n1560(net661_c1,net661);
INTERCONNECT DFFT_315__FPB_n1495_DFFT_316__FPB_n1496(net662_c1,net662);
INTERCONNECT DFFT_299__FPB_n1479_DFFT_300__FPB_n1480(net663_c1,net663);
INTERCONNECT DFFT_219__FPB_n1399_DFFT_220__FPB_n1400(net664_c1,net664);
INTERCONNECT DFFT_459__FPB_n1639_XOR2T_134_R0(net665_c1,net665);
INTERCONNECT DFFT_307__FPB_n1487_AND2T_99_n100(net666_c1,net666);
INTERCONNECT DFFT_500__FPB_n1680_Split_HOLD_1674(net667_c1,net667);
INTERCONNECT DFFT_492__FPB_n1672_DFFT_493__FPB_n1673(net668_c1,net668);
INTERCONNECT DFFT_484__FPB_n1664_DFFT_485__FPB_n1665(net669_c1,net669);
INTERCONNECT DFFT_468__FPB_n1648_DFFT_469__FPB_n1649(net670_c1,net670);
INTERCONNECT DFFT_412__FPB_n1592_DFFT_413__FPB_n1593(net671_c1,net671);
INTERCONNECT DFFT_404__FPB_n1584_DFFT_405__FPB_n1585(net672_c1,net672);
INTERCONNECT DFFT_388__FPB_n1568_DFFT_389__FPB_n1569(net673_c1,net673);
INTERCONNECT DFFT_316__FPB_n1496_DFFT_317__FPB_n1497(net674_c1,net674);
INTERCONNECT DFFT_476__FPB_n1656_AND2T_135_n136(net675_c1,net675);
INTERCONNECT DFFT_396__FPB_n1576_AND2T_123_n124(net676_c1,net676);
INTERCONNECT DFFT_308__FPB_n1488_XOR2T_100_n101(net677_c1,net677);
INTERCONNECT DFFT_501__FPB_n1681_DFFT_502__FPB_n1682(net678_c1,net678);
INTERCONNECT DFFT_493__FPB_n1673_DFFT_494__FPB_n1674(net679_c1,net679);
INTERCONNECT DFFT_485__FPB_n1665_DFFT_486__FPB_n1666(net680_c1,net680);
INTERCONNECT DFFT_477__FPB_n1657_DFFT_478__FPB_n1658(net681_c1,net681);
INTERCONNECT DFFT_469__FPB_n1649_DFFT_470__FPB_n1650(net682_c1,net682);
INTERCONNECT DFFT_413__FPB_n1593_DFFT_414__FPB_n1594(net683_c1,net683);
INTERCONNECT DFFT_405__FPB_n1585_DFFT_406__FPB_n1586(net684_c1,net684);
INTERCONNECT DFFT_397__FPB_n1577_Split_HOLD_1680(net685_c1,net685);
INTERCONNECT DFFT_389__FPB_n1569_DFFT_390__FPB_n1570(net686_c1,net686);
INTERCONNECT DFFT_317__FPB_n1497_DFFT_318__FPB_n1498(net687_c1,net687);
INTERCONNECT DFFT_309__FPB_n1489_DFFT_310__FPB_n1490(net688_c1,net688);
INTERCONNECT DFFT_510__FPB_n1690_DFFT_511_Q3(net689_c1,net689);
INTERCONNECT DFFT_502__FPB_n1682_DFFT_503__FPB_n1683(net690_c1,net690);
INTERCONNECT DFFT_494__FPB_n1674_DFFT_495__FPB_n1675(net691_c1,net691);
INTERCONNECT DFFT_486__FPB_n1666_DFFT_487__FPB_n1667(net692_c1,net692);
INTERCONNECT DFFT_478__FPB_n1658_DFFT_479__FPB_n1659(net693_c1,net693);
INTERCONNECT DFFT_406__FPB_n1586_DFFT_407__FPB_n1587(net694_c1,net694);
INTERCONNECT DFFT_398__FPB_n1578_DFFT_399__FPB_n1579(net695_c1,net695);
INTERCONNECT DFFT_318__FPB_n1498_DFFT_319__FPB_n1499(net696_c1,net696);
INTERCONNECT DFFT_414__FPB_n1594_OR2T_125_n126(net697_c1,net697);
INTERCONNECT DFFT_503__FPB_n1683_DFFT_504__FPB_n1684(net698_c1,net698);
INTERCONNECT DFFT_487__FPB_n1667_DFFT_488__FPB_n1668(net699_c1,net699);
INTERCONNECT DFFT_479__FPB_n1659_DFFT_480__FPB_n1660(net700_c1,net700);
INTERCONNECT DFFT_415__FPB_n1595_DFFT_416__FPB_n1596(net701_c1,net701);
INTERCONNECT DFFT_407__FPB_n1587_DFFT_408__FPB_n1588(net702_c1,net702);
INTERCONNECT DFFT_319__FPB_n1499_DFFT_320__FPB_n1500(net703_c1,net703);
INTERCONNECT DFFT_495__FPB_n1675_AND2T_141_n142(net704_c1,net704);
INTERCONNECT DFFT_399__FPB_n1579_AND2T_124_n125(net705_c1,net705);
INTERCONNECT DFFT_512__FPB_n1692_DFFT_513__FPB_n1693(net706_c1,net706);
INTERCONNECT DFFT_504__FPB_n1684_DFFT_505__FPB_n1685(net707_c1,net707);
INTERCONNECT DFFT_496__FPB_n1676_DFFT_497__FPB_n1677(net708_c1,net708);
INTERCONNECT DFFT_488__FPB_n1668_DFFT_489__FPB_n1669(net709_c1,net709);
INTERCONNECT DFFT_416__FPB_n1596_DFFT_417__FPB_n1597(net710_c1,net710);
INTERCONNECT DFFT_408__FPB_n1588_DFFT_409__FPB_n1589(net711_c1,net711);
INTERCONNECT DFFT_513__FPB_n1693_Split_HOLD_1671(net712_c1,net712);
INTERCONNECT DFFT_505__FPB_n1685_DFFT_506__FPB_n1686(net713_c1,net713);
INTERCONNECT DFFT_497__FPB_n1677_DFFT_498__FPB_n1678(net714_c1,net714);
INTERCONNECT DFFT_489__FPB_n1669_DFFT_490__FPB_n1670(net715_c1,net715);
INTERCONNECT DFFT_417__FPB_n1597_DFFT_418__FPB_n1598(net716_c1,net716);
INTERCONNECT DFFT_409__FPB_n1589_DFFT_410__FPB_n1590(net717_c1,net717);
INTERCONNECT DFFT_514__FPB_n1694_DFFT_515__FPB_n1695(net718_c1,net718);
INTERCONNECT DFFT_506__FPB_n1686_DFFT_507__FPB_n1687(net719_c1,net719);
INTERCONNECT DFFT_498__FPB_n1678_DFFT_499__FPB_n1679(net720_c1,net720);
INTERCONNECT DFFT_418__FPB_n1598_DFFT_419__FPB_n1599(net721_c1,net721);
INTERCONNECT DFFT_515__FPB_n1695_DFFT_516__FPB_n1696(net722_c1,net722);
INTERCONNECT DFFT_507__FPB_n1687_DFFT_508__FPB_n1688(net723_c1,net723);
INTERCONNECT DFFT_499__FPB_n1679_DFFT_500__FPB_n1680(net724_c1,net724);
INTERCONNECT DFFT_419__FPB_n1599_DFFT_420__FPB_n1600(net725_c1,net725);
INTERCONNECT DFFT_516__FPB_n1696_DFFT_517__FPB_n1697(net726_c1,net726);
INTERCONNECT DFFT_508__FPB_n1688_DFFT_509__FPB_n1689(net727_c1,net727);
INTERCONNECT DFFT_517__FPB_n1697_DFFT_518__FPB_n1698(net728_c1,net728);
INTERCONNECT DFFT_509__FPB_n1689_DFFT_510__FPB_n1690(net729_c1,net729);
INTERCONNECT DFFT_518__FPB_n1698_DFFT_519__FPB_n1699(net730_c1,net730);
INTERCONNECT DFFT_519__FPB_n1699_DFFT_520__FPB_n1700(net731_c1,net731);
INTERCONNECT DFFT_142__FPB_n143_Split_626_n1806(net732_c1,net732);
INTERCONNECT DFFT_143__FPB_n144_Split_629_n1809(net733_c1,net733);
INTERCONNECT DFFT_144__FPB_n145_Split_632_n1812(net734_c1,net734);
INTERCONNECT DFFT_145__FPB_n146_Split_635_n1815(net735_c1,net735);
INTERCONNECT DFFT_146__FPB_n147_Split_638_n1818(net736_c1,net736);
INTERCONNECT DFFT_147__FPB_n148_Split_641_n1821(net737_c1,net737);
INTERCONNECT SplitCLK_0_1547_SplitCLK_0_785(net738_c1,net738);
INTERCONNECT SplitCLK_0_1547_SplitCLK_2_1046(net739_c1,net739);
INTERCONNECT SplitCLK_2_1546_DFFT_518__FPB_n1698(net740_c1,net740);
INTERCONNECT SplitCLK_2_1545_DFFT_198__FPB_n1378(net741_c1,net741);
INTERCONNECT SplitCLK_4_1544_DFFT_278__FPB_n1458(net742_c1,net742);
INTERCONNECT SplitCLK_4_1543_DFFT_286__FPB_n1466(net743_c1,net743);
INTERCONNECT SplitCLK_2_1542_DFFT_294__FPB_n1474(net744_c1,net744);
INTERCONNECT SplitCLK_2_1541_DFFT_358__FPB_n1538(net745_c1,net745);
INTERCONNECT SplitCLK_4_1540_DFFT_366__FPB_n1546(net746_c1,net746);
INTERCONNECT SplitCLK_2_1539_DFFT_374__FPB_n1554(net747_c1,net747);
INTERCONNECT SplitCLK_2_1538_DFFT_382__FPB_n1562(net748_c1,net748);
INTERCONNECT SplitCLK_2_1537_DFFT_390__FPB_n1570(net749_c1,net749);
INTERCONNECT SplitCLK_2_1536_DFFT_438__FPB_n1618(net750_c1,net750);
INTERCONNECT SplitCLK_4_1535_DFFT_446__FPB_n1626(net751_c1,net751);
INTERCONNECT SplitCLK_4_1534_DFFT_454__FPB_n1634(net752_c1,net752);
INTERCONNECT SplitCLK_4_1533_DFFT_462__FPB_n1642(net753_c1,net753);
INTERCONNECT SplitCLK_4_1532_DFFT_526__FPB_n1706(net754_c1,net754);
INTERCONNECT SplitCLK_2_1531_DFFT_534__FPB_n1714(net755_c1,net755);
INTERCONNECT SplitCLK_4_1530_DFFT_509__FPB_n1689(net756_c1,net756);
INTERCONNECT SplitCLK_2_1529_DFFT_517__FPB_n1697(net757_c1,net757);
INTERCONNECT SplitCLK_2_1528_DFFT_197__FPB_n1377(net758_c1,net758);
INTERCONNECT SplitCLK_2_1527_DFFT_269__FPB_n1449(net759_c1,net759);
INTERCONNECT SplitCLK_2_1526_DFFT_277__FPB_n1457(net760_c1,net760);
INTERCONNECT SplitCLK_4_1525_DFFT_285__FPB_n1465(net761_c1,net761);
INTERCONNECT SplitCLK_4_1524_DFFT_293__FPB_n1473(net762_c1,net762);
INTERCONNECT SplitCLK_4_1523_DFFT_349__FPB_n1529(net763_c1,net763);
INTERCONNECT SplitCLK_4_1522_DFFT_357__FPB_n1537(net764_c1,net764);
INTERCONNECT SplitCLK_2_1521_DFFT_365__FPB_n1545(net765_c1,net765);
INTERCONNECT SplitCLK_2_1520_DFFT_373__FPB_n1553(net766_c1,net766);
INTERCONNECT SplitCLK_2_1519_DFFT_381__FPB_n1561(net767_c1,net767);
INTERCONNECT SplitCLK_2_1518_DFFT_429__FPB_n1609(net768_c1,net768);
INTERCONNECT SplitCLK_2_1517_DFFT_437__FPB_n1617(net769_c1,net769);
INTERCONNECT SplitCLK_2_1516_DFFT_445__FPB_n1625(net770_c1,net770);
INTERCONNECT SplitCLK_2_1515_DFFT_453__FPB_n1633(net771_c1,net771);
INTERCONNECT SplitCLK_2_1514_DFFT_525__FPB_n1705(net772_c1,net772);
INTERCONNECT SplitCLK_4_1513_DFFT_533__FPB_n1713(net773_c1,net773);
INTERCONNECT SplitCLK_2_1512_DFFT_508__FPB_n1688(net774_c1,net774);
INTERCONNECT SplitCLK_2_1511_DFFT_516__FPB_n1696(net775_c1,net775);
INTERCONNECT SplitCLK_4_1510_DFFT_196__FPB_n1376(net776_c1,net776);
INTERCONNECT SplitCLK_4_1509_DFFT_268__FPB_n1448(net777_c1,net777);
INTERCONNECT SplitCLK_4_1508_DFFT_276__FPB_n1456(net778_c1,net778);
INTERCONNECT SplitCLK_2_1507_DFFT_284__FPB_n1464(net779_c1,net779);
INTERCONNECT SplitCLK_2_1506_DFFT_292__FPB_n1472(net780_c1,net780);
INTERCONNECT SplitCLK_4_1505_DFFT_348__FPB_n1528(net781_c1,net781);
INTERCONNECT SplitCLK_2_1504_DFFT_356__FPB_n1536(net782_c1,net782);
INTERCONNECT SplitCLK_4_1503_DFFT_364__FPB_n1544(net783_c1,net783);
INTERCONNECT SplitCLK_4_1502_DFFT_372__FPB_n1552(net784_c1,net784);
INTERCONNECT SplitCLK_4_1501_DFFT_380__FPB_n1560(net785_c1,net785);
INTERCONNECT SplitCLK_4_1500_DFFT_428__FPB_n1608(net786_c1,net786);
INTERCONNECT SplitCLK_4_1499_DFFT_436__FPB_n1616(net787_c1,net787);
INTERCONNECT SplitCLK_4_1498_DFFT_444__FPB_n1624(net788_c1,net788);
INTERCONNECT SplitCLK_4_1497_DFFT_452__FPB_n1632(net789_c1,net789);
INTERCONNECT SplitCLK_2_1496_DFFT_460__FPB_n1640(net790_c1,net790);
INTERCONNECT SplitCLK_4_1495_DFFT_524__FPB_n1704(net791_c1,net791);
INTERCONNECT SplitCLK_2_1494_DFFT_532__FPB_n1712(net792_c1,net792);
INTERCONNECT SplitCLK_4_1493_DFFT_419__FPB_n1599(net793_c1,net793);
INTERCONNECT SplitCLK_4_1492_DFFT_507__FPB_n1687(net794_c1,net794);
INTERCONNECT SplitCLK_4_1491_DFFT_515__FPB_n1695(net795_c1,net795);
INTERCONNECT SplitCLK_2_1490_DFFT_179__FPB_n1359(net796_c1,net796);
INTERCONNECT SplitCLK_2_1489_DFFT_187__FPB_n1367(net797_c1,net797);
INTERCONNECT SplitCLK_2_1488_DFFT_195__FPB_n1375(net798_c1,net798);
INTERCONNECT SplitCLK_4_1487_DFFT_259__FPB_n1439(net799_c1,net799);
INTERCONNECT SplitCLK_4_1486_DFFT_267__FPB_n1447(net800_c1,net800);
INTERCONNECT SplitCLK_2_1485_DFFT_275__FPB_n1455(net801_c1,net801);
INTERCONNECT SplitCLK_2_1484_DFFT_283__FPB_n1463(net802_c1,net802);
INTERCONNECT SplitCLK_4_1483_DFFT_291__FPB_n1471(net803_c1,net803);
INTERCONNECT SplitCLK_2_1482_DFFT_339__FPB_n1519(net804_c1,net804);
INTERCONNECT SplitCLK_2_1481_DFFT_347__FPB_n1527(net805_c1,net805);
INTERCONNECT SplitCLK_4_1480_DFFT_355__FPB_n1535(net806_c1,net806);
INTERCONNECT SplitCLK_2_1479_DFFT_363__FPB_n1543(net807_c1,net807);
INTERCONNECT SplitCLK_2_1478_DFFT_371__FPB_n1551(net808_c1,net808);
INTERCONNECT SplitCLK_2_1477_DFFT_427__FPB_n1607(net809_c1,net809);
INTERCONNECT SplitCLK_2_1476_DFFT_435__FPB_n1615(net810_c1,net810);
INTERCONNECT SplitCLK_2_1475_DFFT_443__FPB_n1623(net811_c1,net811);
INTERCONNECT SplitCLK_2_1474_DFFT_451__FPB_n1631(net812_c1,net812);
INTERCONNECT SplitCLK_2_1473_DFFT_523__FPB_n1703(net813_c1,net813);
INTERCONNECT SplitCLK_4_1472_DFFT_531__FPB_n1711(net814_c1,net814);
INTERCONNECT SplitCLK_4_1471_NOTT_139_n140(net815_c1,net815);
INTERCONNECT SplitCLK_4_1470_NOTT_138_n139(net816_c1,net816);
INTERCONNECT SplitCLK_2_1469_NOTT_137_n138(net817_c1,net817);
INTERCONNECT SplitCLK_2_1468_NOTT_136_n137(net818_c1,net818);
INTERCONNECT SplitCLK_2_1467_NOTT_107_n108(net819_c1,net819);
INTERCONNECT SplitCLK_4_1466_NOTT_104_n105(net820_c1,net820);
INTERCONNECT SplitCLK_4_1465_NOTT_110_n111(net821_c1,net821);
INTERCONNECT SplitCLK_2_1464_NOTT_101_n102(net822_c1,net822);
INTERCONNECT SplitCLK_2_1463_DFFT_418__FPB_n1598(net823_c1,net823);
INTERCONNECT SplitCLK_4_1462_DFFT_506__FPB_n1686(net824_c1,net824);
INTERCONNECT SplitCLK_2_1461_DFFT_514__FPB_n1694(net825_c1,net825);
INTERCONNECT SplitCLK_2_1460_DFFT_178__FPB_n1358(net826_c1,net826);
INTERCONNECT SplitCLK_4_1459_DFFT_186__FPB_n1366(net827_c1,net827);
INTERCONNECT SplitCLK_2_1458_DFFT_194__FPB_n1374(net828_c1,net828);
INTERCONNECT SplitCLK_2_1457_DFFT_258__FPB_n1438(net829_c1,net829);
INTERCONNECT SplitCLK_2_1456_DFFT_266__FPB_n1446(net830_c1,net830);
INTERCONNECT SplitCLK_2_1455_DFFT_274__FPB_n1454(net831_c1,net831);
INTERCONNECT SplitCLK_2_1454_DFFT_282__FPB_n1462(net832_c1,net832);
INTERCONNECT SplitCLK_2_1453_DFFT_290__FPB_n1470(net833_c1,net833);
INTERCONNECT SplitCLK_4_1452_DFFT_338__FPB_n1518(net834_c1,net834);
INTERCONNECT SplitCLK_4_1451_DFFT_346__FPB_n1526(net835_c1,net835);
INTERCONNECT SplitCLK_2_1450_DFFT_354__FPB_n1534(net836_c1,net836);
INTERCONNECT SplitCLK_2_1449_DFFT_362__FPB_n1542(net837_c1,net837);
INTERCONNECT SplitCLK_4_1448_DFFT_370__FPB_n1550(net838_c1,net838);
INTERCONNECT SplitCLK_4_1447_DFFT_426__FPB_n1606(net839_c1,net839);
INTERCONNECT SplitCLK_2_1446_DFFT_434__FPB_n1614(net840_c1,net840);
INTERCONNECT SplitCLK_4_1445_DFFT_442__FPB_n1622(net841_c1,net841);
INTERCONNECT SplitCLK_4_1444_DFFT_450__FPB_n1630(net842_c1,net842);
INTERCONNECT SplitCLK_2_1443_DFFT_530__FPB_n1710(net843_c1,net843);
INTERCONNECT SplitCLK_4_1442_DFFT_409__FPB_n1589(net844_c1,net844);
INTERCONNECT SplitCLK_4_1441_DFFT_417__FPB_n1597(net845_c1,net845);
INTERCONNECT SplitCLK_2_1440_DFFT_505__FPB_n1685(net846_c1,net846);
INTERCONNECT SplitCLK_4_1439_DFFT_513__FPB_n1693(net847_c1,net847);
INTERCONNECT SplitCLK_2_1438_DFFT_169__FPB_n1349(net848_c1,net848);
INTERCONNECT SplitCLK_2_1437_DFFT_177__FPB_n1357(net849_c1,net849);
INTERCONNECT SplitCLK_2_1436_DFFT_185__FPB_n1365(net850_c1,net850);
INTERCONNECT SplitCLK_4_1435_DFFT_193__FPB_n1373(net851_c1,net851);
INTERCONNECT SplitCLK_2_1434_DFFT_249__FPB_n1429(net852_c1,net852);
INTERCONNECT SplitCLK_4_1433_DFFT_257__FPB_n1437(net853_c1,net853);
INTERCONNECT SplitCLK_4_1432_DFFT_265__FPB_n1445(net854_c1,net854);
INTERCONNECT SplitCLK_2_1431_DFFT_273__FPB_n1453(net855_c1,net855);
INTERCONNECT SplitCLK_4_1430_DFFT_281__FPB_n1461(net856_c1,net856);
INTERCONNECT SplitCLK_2_1429_DFFT_329__FPB_n1509(net857_c1,net857);
INTERCONNECT SplitCLK_2_1428_DFFT_337__FPB_n1517(net858_c1,net858);
INTERCONNECT SplitCLK_4_1427_DFFT_345__FPB_n1525(net859_c1,net859);
INTERCONNECT SplitCLK_4_1426_DFFT_361__FPB_n1541(net860_c1,net860);
INTERCONNECT SplitCLK_2_1425_DFFT_425__FPB_n1605(net861_c1,net861);
INTERCONNECT SplitCLK_2_1424_DFFT_433__FPB_n1613(net862_c1,net862);
INTERCONNECT SplitCLK_2_1423_DFFT_441__FPB_n1621(net863_c1,net863);
INTERCONNECT SplitCLK_2_1422_DFFT_521__FPB_n1701(net864_c1,net864);
INTERCONNECT SplitCLK_2_1421_DFFT_147__FPB_n148(net865_c1,net865);
INTERCONNECT SplitCLK_4_1420_DFFT_146__FPB_n147(net866_c1,net866);
INTERCONNECT SplitCLK_4_1419_DFFT_408__FPB_n1588(net867_c1,net867);
INTERCONNECT SplitCLK_2_1418_DFFT_416__FPB_n1596(net868_c1,net868);
INTERCONNECT SplitCLK_4_1417_DFFT_504__FPB_n1684(net869_c1,net869);
INTERCONNECT SplitCLK_2_1416_DFFT_512__FPB_n1692(net870_c1,net870);
INTERCONNECT SplitCLK_4_1415_DFFT_168__FPB_n1348(net871_c1,net871);
INTERCONNECT SplitCLK_2_1414_DFFT_176__FPB_n1356(net872_c1,net872);
INTERCONNECT SplitCLK_4_1413_DFFT_184__FPB_n1364(net873_c1,net873);
INTERCONNECT SplitCLK_4_1412_DFFT_248__FPB_n1428(net874_c1,net874);
INTERCONNECT SplitCLK_4_1411_DFFT_256__FPB_n1436(net875_c1,net875);
INTERCONNECT SplitCLK_4_1410_DFFT_264__FPB_n1444(net876_c1,net876);
INTERCONNECT SplitCLK_4_1409_DFFT_272__FPB_n1452(net877_c1,net877);
INTERCONNECT SplitCLK_4_1408_DFFT_280__FPB_n1460(net878_c1,net878);
INTERCONNECT SplitCLK_4_1407_DFFT_328__FPB_n1508(net879_c1,net879);
INTERCONNECT SplitCLK_4_1406_DFFT_336__FPB_n1516(net880_c1,net880);
INTERCONNECT SplitCLK_2_1405_DFFT_344__FPB_n1524(net881_c1,net881);
INTERCONNECT SplitCLK_2_1404_DFFT_352__FPB_n1532(net882_c1,net882);
INTERCONNECT SplitCLK_2_1403_DFFT_360__FPB_n1540(net883_c1,net883);
INTERCONNECT SplitCLK_4_1402_DFFT_424__FPB_n1604(net884_c1,net884);
INTERCONNECT SplitCLK_4_1401_DFFT_432__FPB_n1612(net885_c1,net885);
INTERCONNECT SplitCLK_4_1400_DFFT_440__FPB_n1620(net886_c1,net886);
INTERCONNECT SplitCLK_2_1399_DFFT_520__FPB_n1700(net887_c1,net887);
INTERCONNECT SplitCLK_2_1398_DFFT_145__FPB_n146(net888_c1,net888);
INTERCONNECT SplitCLK_4_1397_DFFT_144__FPB_n145(net889_c1,net889);
INTERCONNECT SplitCLK_4_1396_DFFT_319__FPB_n1499(net890_c1,net890);
INTERCONNECT SplitCLK_2_1395_DFFT_407__FPB_n1587(net891_c1,net891);
INTERCONNECT SplitCLK_2_1394_DFFT_415__FPB_n1595(net892_c1,net892);
INTERCONNECT SplitCLK_2_1393_DFFT_503__FPB_n1683(net893_c1,net893);
INTERCONNECT SplitCLK_4_1392_DFFT_159__FPB_n1339(net894_c1,net894);
INTERCONNECT SplitCLK_2_1391_DFFT_167__FPB_n1347(net895_c1,net895);
INTERCONNECT SplitCLK_4_1390_DFFT_175__FPB_n1355(net896_c1,net896);
INTERCONNECT SplitCLK_2_1389_DFFT_183__FPB_n1363(net897_c1,net897);
INTERCONNECT SplitCLK_4_1388_DFFT_191__FPB_n1371(net898_c1,net898);
INTERCONNECT SplitCLK_4_1387_DFFT_239__FPB_n1419(net899_c1,net899);
INTERCONNECT SplitCLK_4_1386_DFFT_247__FPB_n1427(net900_c1,net900);
INTERCONNECT SplitCLK_2_1385_DFFT_255__FPB_n1435(net901_c1,net901);
INTERCONNECT SplitCLK_2_1384_DFFT_263__FPB_n1443(net902_c1,net902);
INTERCONNECT SplitCLK_2_1383_DFFT_271__FPB_n1451(net903_c1,net903);
INTERCONNECT SplitCLK_2_1382_DFFT_327__FPB_n1507(net904_c1,net904);
INTERCONNECT SplitCLK_2_1381_DFFT_335__FPB_n1515(net905_c1,net905);
INTERCONNECT SplitCLK_2_1380_DFFT_343__FPB_n1523(net906_c1,net906);
INTERCONNECT SplitCLK_4_1379_DFFT_351__FPB_n1531(net907_c1,net907);
INTERCONNECT SplitCLK_4_1378_DFFT_423__FPB_n1603(net908_c1,net908);
INTERCONNECT SplitCLK_4_1377_DFFT_431__FPB_n1611(net909_c1,net909);
INTERCONNECT SplitCLK_4_1376_DFFT_142__FPB_n143(net910_c1,net910);
INTERCONNECT SplitCLK_2_1375_DFFT_318__FPB_n1498(net911_c1,net911);
INTERCONNECT SplitCLK_4_1374_DFFT_406__FPB_n1586(net912_c1,net912);
INTERCONNECT SplitCLK_2_1373_DFFT_414__FPB_n1594(net913_c1,net913);
INTERCONNECT SplitCLK_4_1372_DFFT_502__FPB_n1682(net914_c1,net914);
INTERCONNECT SplitCLK_4_1371_DFFT_510__FPB_n1690(net915_c1,net915);
INTERCONNECT SplitCLK_4_1370_DFFT_158__FPB_n1338(net916_c1,net916);
INTERCONNECT SplitCLK_4_1369_DFFT_166__FPB_n1346(net917_c1,net917);
INTERCONNECT SplitCLK_2_1368_DFFT_174__FPB_n1354(net918_c1,net918);
INTERCONNECT SplitCLK_4_1367_DFFT_182__FPB_n1362(net919_c1,net919);
INTERCONNECT SplitCLK_4_1366_DFFT_190__FPB_n1370(net920_c1,net920);
INTERCONNECT SplitCLK_2_1365_DFFT_238__FPB_n1418(net921_c1,net921);
INTERCONNECT SplitCLK_2_1364_DFFT_246__FPB_n1426(net922_c1,net922);
INTERCONNECT SplitCLK_4_1363_DFFT_254__FPB_n1434(net923_c1,net923);
INTERCONNECT SplitCLK_2_1362_DFFT_262__FPB_n1442(net924_c1,net924);
INTERCONNECT SplitCLK_4_1361_DFFT_270__FPB_n1450(net925_c1,net925);
INTERCONNECT SplitCLK_2_1360_DFFT_326__FPB_n1506(net926_c1,net926);
INTERCONNECT SplitCLK_2_1359_DFFT_334__FPB_n1514(net927_c1,net927);
INTERCONNECT SplitCLK_4_1358_DFFT_342__FPB_n1522(net928_c1,net928);
INTERCONNECT SplitCLK_2_1357_DFFT_350__FPB_n1530(net929_c1,net929);
INTERCONNECT SplitCLK_4_1356_DFFT_422__FPB_n1602(net930_c1,net930);
INTERCONNECT SplitCLK_4_1355_DFFT_430__FPB_n1610(net931_c1,net931);
INTERCONNECT SplitCLK_2_1354_DFFT_309__FPB_n1489(net932_c1,net932);
INTERCONNECT SplitCLK_4_1353_DFFT_317__FPB_n1497(net933_c1,net933);
INTERCONNECT SplitCLK_2_1352_DFFT_405__FPB_n1585(net934_c1,net934);
INTERCONNECT SplitCLK_4_1351_DFFT_413__FPB_n1593(net935_c1,net935);
INTERCONNECT SplitCLK_4_1350_DFFT_501__FPB_n1681(net936_c1,net936);
INTERCONNECT SplitCLK_4_1349_DFFT_149__FPB_n1329(net937_c1,net937);
INTERCONNECT SplitCLK_2_1348_DFFT_157__FPB_n1337(net938_c1,net938);
INTERCONNECT SplitCLK_4_1347_DFFT_165__FPB_n1345(net939_c1,net939);
INTERCONNECT SplitCLK_2_1346_DFFT_173__FPB_n1353(net940_c1,net940);
INTERCONNECT SplitCLK_2_1345_DFFT_181__FPB_n1361(net941_c1,net941);
INTERCONNECT SplitCLK_2_1344_DFFT_229__FPB_n1409(net942_c1,net942);
INTERCONNECT SplitCLK_2_1343_DFFT_237__FPB_n1417(net943_c1,net943);
INTERCONNECT SplitCLK_2_1342_DFFT_245__FPB_n1425(net944_c1,net944);
INTERCONNECT SplitCLK_4_1341_DFFT_253__FPB_n1433(net945_c1,net945);
INTERCONNECT SplitCLK_4_1340_DFFT_261__FPB_n1441(net946_c1,net946);
INTERCONNECT SplitCLK_2_1339_DFFT_325__FPB_n1505(net947_c1,net947);
INTERCONNECT SplitCLK_4_1338_DFFT_333__FPB_n1513(net948_c1,net948);
INTERCONNECT SplitCLK_2_1337_DFFT_341__FPB_n1521(net949_c1,net949);
INTERCONNECT SplitCLK_2_1336_DFFT_421__FPB_n1601(net950_c1,net950);
INTERCONNECT SplitCLK_4_1335_DFFT_308__FPB_n1488(net951_c1,net951);
INTERCONNECT SplitCLK_4_1334_DFFT_316__FPB_n1496(net952_c1,net952);
INTERCONNECT SplitCLK_4_1333_DFFT_404__FPB_n1584(net953_c1,net953);
INTERCONNECT SplitCLK_4_1332_DFFT_412__FPB_n1592(net954_c1,net954);
INTERCONNECT SplitCLK_2_1331_DFFT_500__FPB_n1680(net955_c1,net955);
INTERCONNECT SplitCLK_4_1330_DFFT_148__FPB_n1328(net956_c1,net956);
INTERCONNECT SplitCLK_2_1329_DFFT_156__FPB_n1336(net957_c1,net957);
INTERCONNECT SplitCLK_2_1328_DFFT_164__FPB_n1344(net958_c1,net958);
INTERCONNECT SplitCLK_4_1327_DFFT_172__FPB_n1352(net959_c1,net959);
INTERCONNECT SplitCLK_4_1326_DFFT_180__FPB_n1360(net960_c1,net960);
INTERCONNECT SplitCLK_4_1325_DFFT_228__FPB_n1408(net961_c1,net961);
INTERCONNECT SplitCLK_2_1324_DFFT_244__FPB_n1424(net962_c1,net962);
INTERCONNECT SplitCLK_2_1323_DFFT_252__FPB_n1432(net963_c1,net963);
INTERCONNECT SplitCLK_2_1322_DFFT_260__FPB_n1440(net964_c1,net964);
INTERCONNECT SplitCLK_2_1321_DFFT_324__FPB_n1504(net965_c1,net965);
INTERCONNECT SplitCLK_2_1320_DFFT_332__FPB_n1512(net966_c1,net966);
INTERCONNECT SplitCLK_2_1319_DFFT_340__FPB_n1520(net967_c1,net967);
INTERCONNECT SplitCLK_2_1318_DFFT_420__FPB_n1600(net968_c1,net968);
INTERCONNECT SplitCLK_2_1317_DFFT_219__FPB_n1399(net969_c1,net969);
INTERCONNECT SplitCLK_4_1316_DFFT_307__FPB_n1487(net970_c1,net970);
INTERCONNECT SplitCLK_2_1315_DFFT_315__FPB_n1495(net971_c1,net971);
INTERCONNECT SplitCLK_2_1314_DFFT_403__FPB_n1583(net972_c1,net972);
INTERCONNECT SplitCLK_4_1313_DFFT_411__FPB_n1591(net973_c1,net973);
INTERCONNECT SplitCLK_2_1312_DFFT_155__FPB_n1335(net974_c1,net974);
INTERCONNECT SplitCLK_4_1311_DFFT_163__FPB_n1343(net975_c1,net975);
INTERCONNECT SplitCLK_2_1310_DFFT_171__FPB_n1351(net976_c1,net976);
INTERCONNECT SplitCLK_2_1309_DFFT_227__FPB_n1407(net977_c1,net977);
INTERCONNECT SplitCLK_4_1308_DFFT_235__FPB_n1415(net978_c1,net978);
INTERCONNECT SplitCLK_4_1307_DFFT_243__FPB_n1423(net979_c1,net979);
INTERCONNECT SplitCLK_2_1306_DFFT_251__FPB_n1431(net980_c1,net980);
INTERCONNECT SplitCLK_4_1305_DFFT_323__FPB_n1503(net981_c1,net981);
INTERCONNECT SplitCLK_2_1304_DFFT_331__FPB_n1511(net982_c1,net982);
INTERCONNECT SplitCLK_4_1303_DFFT_218__FPB_n1398(net983_c1,net983);
INTERCONNECT SplitCLK_4_1302_DFFT_306__FPB_n1486(net984_c1,net984);
INTERCONNECT SplitCLK_4_1301_DFFT_314__FPB_n1494(net985_c1,net985);
INTERCONNECT SplitCLK_2_1300_DFFT_402__FPB_n1582(net986_c1,net986);
INTERCONNECT SplitCLK_2_1299_DFFT_410__FPB_n1590(net987_c1,net987);
INTERCONNECT SplitCLK_2_1298_DFFT_154__FPB_n1334(net988_c1,net988);
INTERCONNECT SplitCLK_2_1297_DFFT_162__FPB_n1342(net989_c1,net989);
INTERCONNECT SplitCLK_4_1296_DFFT_170__FPB_n1350(net990_c1,net990);
INTERCONNECT SplitCLK_4_1295_DFFT_226__FPB_n1406(net991_c1,net991);
INTERCONNECT SplitCLK_2_1294_DFFT_234__FPB_n1414(net992_c1,net992);
INTERCONNECT SplitCLK_2_1293_DFFT_242__FPB_n1422(net993_c1,net993);
INTERCONNECT SplitCLK_4_1292_DFFT_250__FPB_n1430(net994_c1,net994);
INTERCONNECT SplitCLK_4_1291_DFFT_322__FPB_n1502(net995_c1,net995);
INTERCONNECT SplitCLK_4_1290_DFFT_330__FPB_n1510(net996_c1,net996);
INTERCONNECT SplitCLK_4_1289_AND2T_99_n100(net997_c1,net997);
INTERCONNECT SplitCLK_2_1288_DFFT_209__FPB_n1389(net998_c1,net998);
INTERCONNECT SplitCLK_2_1287_DFFT_217__FPB_n1397(net999_c1,net999);
INTERCONNECT SplitCLK_2_1286_DFFT_305__FPB_n1485(net1000_c1,net1000);
INTERCONNECT SplitCLK_2_1285_DFFT_313__FPB_n1493(net1001_c1,net1001);
INTERCONNECT SplitCLK_2_1284_DFFT_401__FPB_n1581(net1002_c1,net1002);
INTERCONNECT SplitCLK_4_1283_DFFT_153__FPB_n1333(net1003_c1,net1003);
INTERCONNECT SplitCLK_4_1282_DFFT_161__FPB_n1341(net1004_c1,net1004);
INTERCONNECT SplitCLK_4_1281_DFFT_225__FPB_n1405(net1005_c1,net1005);
INTERCONNECT SplitCLK_2_1280_DFFT_233__FPB_n1413(net1006_c1,net1006);
INTERCONNECT SplitCLK_4_1279_DFFT_241__FPB_n1421(net1007_c1,net1007);
INTERCONNECT SplitCLK_2_1278_DFFT_321__FPB_n1501(net1008_c1,net1008);
INTERCONNECT SplitCLK_2_1277_DFFT_208__FPB_n1388(net1009_c1,net1009);
INTERCONNECT SplitCLK_4_1276_DFFT_216__FPB_n1396(net1010_c1,net1010);
INTERCONNECT SplitCLK_2_1275_DFFT_304__FPB_n1484(net1011_c1,net1011);
INTERCONNECT SplitCLK_4_1274_DFFT_312__FPB_n1492(net1012_c1,net1012);
INTERCONNECT SplitCLK_4_1273_DFFT_400__FPB_n1580(net1013_c1,net1013);
INTERCONNECT SplitCLK_2_1272_DFFT_160__FPB_n1340(net1014_c1,net1014);
INTERCONNECT SplitCLK_2_1271_DFFT_224__FPB_n1404(net1015_c1,net1015);
INTERCONNECT SplitCLK_2_1270_DFFT_232__FPB_n1412(net1016_c1,net1016);
INTERCONNECT SplitCLK_2_1269_DFFT_240__FPB_n1420(net1017_c1,net1017);
INTERCONNECT SplitCLK_4_1268_DFFT_320__FPB_n1500(net1018_c1,net1018);
INTERCONNECT SplitCLK_2_1267_DFFT_207__FPB_n1387(net1019_c1,net1019);
INTERCONNECT SplitCLK_4_1266_DFFT_215__FPB_n1395(net1020_c1,net1020);
INTERCONNECT SplitCLK_4_1265_DFFT_303__FPB_n1483(net1021_c1,net1021);
INTERCONNECT SplitCLK_2_1264_DFFT_311__FPB_n1491(net1022_c1,net1022);
INTERCONNECT SplitCLK_2_1263_DFFT_223__FPB_n1403(net1023_c1,net1023);
INTERCONNECT SplitCLK_2_1262_XOR2T_128_n129(net1024_c1,net1024);
INTERCONNECT SplitCLK_2_1261_OR2T_119_n120(net1025_c1,net1025);
INTERCONNECT SplitCLK_2_1260_XOR2T_117_n118(net1026_c1,net1026);
INTERCONNECT SplitCLK_2_1259_OR2T_125_n126(net1027_c1,net1027);
INTERCONNECT SplitCLK_2_1258_OR2T_108_n109(net1028_c1,net1028);
INTERCONNECT SplitCLK_4_1257_OR2T_115_n116(net1029_c1,net1029);
INTERCONNECT SplitCLK_2_1256_XOR2T_122_n123(net1030_c1,net1030);
INTERCONNECT SplitCLK_2_1255_OR2T_130_n131(net1031_c1,net1031);
INTERCONNECT SplitCLK_4_1254_XOR2T_105_n106(net1032_c1,net1032);
INTERCONNECT SplitCLK_2_1253_OR2T_113_n114(net1033_c1,net1033);
INTERCONNECT SplitCLK_2_1252_OR2T_102_n103(net1034_c1,net1034);
INTERCONNECT SplitCLK_2_1251_XOR2T_100_n101(net1035_c1,net1035);
INTERCONNECT SplitCLK_2_1250_DFFT_206__FPB_n1386(net1036_c1,net1036);
INTERCONNECT SplitCLK_2_1249_DFFT_302__FPB_n1482(net1037_c1,net1037);
INTERCONNECT SplitCLK_4_1248_DFFT_310__FPB_n1490(net1038_c1,net1038);
INTERCONNECT SplitCLK_2_1247_DFFT_150__FPB_n1330(net1039_c1,net1039);
INTERCONNECT SplitCLK_4_1246_DFFT_222__FPB_n1402(net1040_c1,net1040);
INTERCONNECT SplitCLK_4_1245_DFFT_230__FPB_n1410(net1041_c1,net1041);
INTERCONNECT SplitCLK_2_1244_NOTT_97_n98(net1042_c1,net1042);
INTERCONNECT SplitCLK_2_1243_NOTT_94_n95(net1043_c1,net1043);
INTERCONNECT SplitCLK_2_1242_NOTT_77_n78(net1044_c1,net1044);
INTERCONNECT SplitCLK_2_1241_NOTT_83_n84(net1045_c1,net1045);
INTERCONNECT SplitCLK_4_1240_NOTT_58_n59(net1046_c1,net1046);
INTERCONNECT SplitCLK_4_1239_NOTT_56_n57(net1047_c1,net1047);
INTERCONNECT SplitCLK_2_1238_NOTT_55_n56(net1048_c1,net1048);
INTERCONNECT SplitCLK_2_1237_NOTT_70_n71(net1049_c1,net1049);
INTERCONNECT SplitCLK_2_1236_NOTT_18_n18(net1050_c1,net1050);
INTERCONNECT SplitCLK_2_1235_NOTT_17_n17(net1051_c1,net1051);
INTERCONNECT SplitCLK_2_1234_NOTT_32_n33(net1052_c1,net1052);
INTERCONNECT SplitCLK_4_1233_NOTT_21_n21(net1053_c1,net1053);
INTERCONNECT SplitCLK_2_1232_NOTT_20_n20(net1054_c1,net1054);
INTERCONNECT SplitCLK_2_1231_DFFT_205__FPB_n1385(net1055_c1,net1055);
INTERCONNECT SplitCLK_2_1230_DFFT_213__FPB_n1393(net1056_c1,net1056);
INTERCONNECT SplitCLK_2_1229_DFFT_301__FPB_n1481(net1057_c1,net1057);
INTERCONNECT SplitCLK_4_1228_DFFT_221__FPB_n1401(net1058_c1,net1058);
INTERCONNECT SplitCLK_2_1227_DFFT_204__FPB_n1384(net1059_c1,net1059);
INTERCONNECT SplitCLK_4_1226_DFFT_212__FPB_n1392(net1060_c1,net1060);
INTERCONNECT SplitCLK_4_1225_DFFT_300__FPB_n1480(net1061_c1,net1061);
INTERCONNECT SplitCLK_4_1224_DFFT_220__FPB_n1400(net1062_c1,net1062);
INTERCONNECT SplitCLK_4_1223_DFFT_499__FPB_n1679(net1063_c1,net1063);
INTERCONNECT SplitCLK_2_1222_DFFT_203__FPB_n1383(net1064_c1,net1064);
INTERCONNECT SplitCLK_2_1221_DFFT_211__FPB_n1391(net1065_c1,net1065);
INTERCONNECT SplitCLK_4_1220_OR2T_98_n99(net1066_c1,net1066);
INTERCONNECT SplitCLK_2_1219_OR2T_96_n97(net1067_c1,net1067);
INTERCONNECT SplitCLK_2_1218_OR2T_86_n87(net1068_c1,net1068);
INTERCONNECT SplitCLK_4_1217_OR2T_68_n69(net1069_c1,net1069);
INTERCONNECT SplitCLK_2_1216_OR2T_84_n85(net1070_c1,net1070);
INTERCONNECT SplitCLK_2_1215_OR2T_90_n91(net1071_c1,net1071);
INTERCONNECT SplitCLK_4_1214_OR2T_73_n74(net1072_c1,net1072);
INTERCONNECT SplitCLK_4_1213_OR2T_81_n82(net1073_c1,net1073);
INTERCONNECT SplitCLK_2_1212_OR2T_48_n49(net1074_c1,net1074);
INTERCONNECT SplitCLK_2_1211_OR2T_64_n65(net1075_c1,net1075);
INTERCONNECT SplitCLK_4_1210_OR2T_80_n81(net1076_c1,net1076);
INTERCONNECT SplitCLK_4_1209_OR2T_63_n64(net1077_c1,net1077);
INTERCONNECT SplitCLK_4_1208_OR2T_71_n72(net1078_c1,net1078);
INTERCONNECT SplitCLK_4_1207_OR2T_39_n40(net1079_c1,net1079);
INTERCONNECT SplitCLK_4_1206_OR2T_46_n47(net1080_c1,net1080);
INTERCONNECT SplitCLK_2_1205_OR2T_37_n38(net1081_c1,net1081);
INTERCONNECT SplitCLK_4_1204_OR2T_45_n46(net1082_c1,net1082);
INTERCONNECT SplitCLK_2_1203_OR2T_36_n37(net1083_c1,net1083);
INTERCONNECT SplitCLK_4_1202_OR2T_52_n53(net1084_c1,net1084);
INTERCONNECT SplitCLK_2_1201_OR2T_60_n61(net1085_c1,net1085);
INTERCONNECT SplitCLK_4_1200_OR2T_51_n52(net1086_c1,net1086);
INTERCONNECT SplitCLK_2_1199_OR2T_34_n35(net1087_c1,net1087);
INTERCONNECT SplitCLK_4_1198_OR2T_26_n26(net1088_c1,net1088);
INTERCONNECT SplitCLK_2_1197_OR2T_41_n42(net1089_c1,net1089);
INTERCONNECT SplitCLK_2_1196_OR2T_25_n25(net1090_c1,net1090);
INTERCONNECT SplitCLK_4_1195_OR2T_40_n41(net1091_c1,net1091);
INTERCONNECT SplitCLK_2_1194_OR2T_31_n32(net1092_c1,net1092);
INTERCONNECT SplitCLK_2_1193_OR2T_30_n31(net1093_c1,net1093);
INTERCONNECT SplitCLK_4_1192_OR2T_22_n22(net1094_c1,net1094);
INTERCONNECT SplitCLK_4_1191_OR2T_127_R2(net1095_c1,net1095);
INTERCONNECT SplitCLK_2_1190_OR2T_133_R1(net1096_c1,net1096);
INTERCONNECT SplitCLK_4_1189_DFFT_498__FPB_n1678(net1097_c1,net1097);
INTERCONNECT SplitCLK_2_1188_DFFT_202__FPB_n1382(net1098_c1,net1098);
INTERCONNECT SplitCLK_4_1187_DFFT_210__FPB_n1390(net1099_c1,net1099);
INTERCONNECT SplitCLK_4_1186_DFFT_489__FPB_n1669(net1100_c1,net1100);
INTERCONNECT SplitCLK_2_1185_DFFT_497__FPB_n1677(net1101_c1,net1101);
INTERCONNECT SplitCLK_4_1184_DFFT_201__FPB_n1381(net1102_c1,net1102);
INTERCONNECT SplitCLK_2_1183_DFFT_488__FPB_n1668(net1103_c1,net1103);
INTERCONNECT SplitCLK_4_1182_DFFT_496__FPB_n1676(net1104_c1,net1104);
INTERCONNECT SplitCLK_4_1181_DFFT_200__FPB_n1380(net1105_c1,net1105);
INTERCONNECT SplitCLK_2_1180_AND2T_88_n89(net1106_c1,net1106);
INTERCONNECT SplitCLK_2_1179_AND2T_87_n88(net1107_c1,net1107);
INTERCONNECT SplitCLK_4_1178_AND2T_95_n96(net1108_c1,net1108);
INTERCONNECT SplitCLK_2_1177_AND2T_78_n79(net1109_c1,net1109);
INTERCONNECT SplitCLK_4_1176_AND2T_85_n86(net1110_c1,net1110);
INTERCONNECT SplitCLK_4_1175_AND2T_69_n70(net1111_c1,net1111);
INTERCONNECT SplitCLK_4_1174_AND2T_76_n77(net1112_c1,net1112);
INTERCONNECT SplitCLK_2_1173_AND2T_92_n93(net1113_c1,net1113);
INTERCONNECT SplitCLK_2_1172_AND2T_67_n68(net1114_c1,net1114);
INTERCONNECT SplitCLK_4_1171_AND2T_75_n76(net1115_c1,net1115);
INTERCONNECT SplitCLK_2_1170_AND2T_59_n60(net1116_c1,net1116);
INTERCONNECT SplitCLK_4_1169_AND2T_66_n67(net1117_c1,net1117);
INTERCONNECT SplitCLK_4_1168_AND2T_82_n83(net1118_c1,net1118);
INTERCONNECT SplitCLK_2_1167_AND2T_57_n58(net1119_c1,net1119);
INTERCONNECT SplitCLK_4_1166_AND2T_49_n50(net1120_c1,net1120);
INTERCONNECT SplitCLK_2_1165_AND2T_38_n39(net1121_c1,net1121);
INTERCONNECT SplitCLK_2_1164_AND2T_54_n55(net1122_c1,net1122);
INTERCONNECT SplitCLK_4_1163_AND2T_53_n54(net1123_c1,net1123);
INTERCONNECT SplitCLK_2_1162_AND2T_61_n62(net1124_c1,net1124);
INTERCONNECT SplitCLK_2_1161_AND2T_29_n30(net1125_c1,net1125);
INTERCONNECT SplitCLK_4_1160_AND2T_28_n28(net1126_c1,net1126);
INTERCONNECT SplitCLK_4_1159_AND2T_35_n36(net1127_c1,net1127);
INTERCONNECT SplitCLK_2_1158_AND2T_43_n44(net1128_c1,net1128);
INTERCONNECT SplitCLK_2_1157_AND2T_19_n19(net1129_c1,net1129);
INTERCONNECT SplitCLK_2_1156_AND2T_27_n27(net1130_c1,net1130);
INTERCONNECT SplitCLK_4_1155_AND2T_42_n43(net1131_c1,net1131);
INTERCONNECT SplitCLK_2_1154_AND2T_50_n51(net1132_c1,net1132);
INTERCONNECT SplitCLK_4_1153_AND2T_33_n34(net1133_c1,net1133);
INTERCONNECT SplitCLK_2_1152_AND2T_24_n24(net1134_c1,net1134);
INTERCONNECT SplitCLK_2_1151_AND2T_23_n23(net1135_c1,net1135);
INTERCONNECT SplitCLK_2_1150_AND2T_120_R3(net1136_c1,net1136);
INTERCONNECT SplitCLK_2_1149_DFFT_399__FPB_n1579(net1137_c1,net1137);
INTERCONNECT SplitCLK_2_1148_DFFT_479__FPB_n1659(net1138_c1,net1138);
INTERCONNECT SplitCLK_4_1147_DFFT_487__FPB_n1667(net1139_c1,net1139);
INTERCONNECT SplitCLK_4_1146_DFFT_495__FPB_n1675(net1140_c1,net1140);
INTERCONNECT SplitCLK_4_1145_DFFT_398__FPB_n1578(net1141_c1,net1141);
INTERCONNECT SplitCLK_4_1144_DFFT_478__FPB_n1658(net1142_c1,net1142);
INTERCONNECT SplitCLK_2_1143_DFFT_486__FPB_n1666(net1143_c1,net1143);
INTERCONNECT SplitCLK_2_1142_DFFT_494__FPB_n1674(net1144_c1,net1144);
INTERCONNECT SplitCLK_2_1141_DFFT_389__FPB_n1569(net1145_c1,net1145);
INTERCONNECT SplitCLK_2_1140_DFFT_397__FPB_n1577(net1146_c1,net1146);
INTERCONNECT SplitCLK_4_1139_DFFT_477__FPB_n1657(net1147_c1,net1147);
INTERCONNECT SplitCLK_4_1138_DFFT_485__FPB_n1665(net1148_c1,net1148);
INTERCONNECT SplitCLK_2_1137_DFFT_493__FPB_n1673(net1149_c1,net1149);
INTERCONNECT SplitCLK_2_1136_DFFT_527_Q2(net1150_c1,net1150);
INTERCONNECT SplitCLK_2_1135_DFFT_540_Q0(net1151_c1,net1151);
INTERCONNECT SplitCLK_2_1134_DFFT_511_Q3(net1152_c1,net1152);
INTERCONNECT SplitCLK_2_1133_DFFT_388__FPB_n1568(net1153_c1,net1153);
INTERCONNECT SplitCLK_4_1132_DFFT_396__FPB_n1576(net1154_c1,net1154);
INTERCONNECT SplitCLK_4_1131_DFFT_468__FPB_n1648(net1155_c1,net1155);
INTERCONNECT SplitCLK_2_1130_DFFT_476__FPB_n1656(net1156_c1,net1156);
INTERCONNECT SplitCLK_2_1129_DFFT_484__FPB_n1664(net1157_c1,net1157);
INTERCONNECT SplitCLK_4_1128_DFFT_492__FPB_n1672(net1158_c1,net1158);
INTERCONNECT SplitCLK_2_1127_DFFT_299__FPB_n1479(net1159_c1,net1159);
INTERCONNECT SplitCLK_2_1126_DFFT_379__FPB_n1559(net1160_c1,net1160);
INTERCONNECT SplitCLK_4_1125_DFFT_387__FPB_n1567(net1161_c1,net1161);
INTERCONNECT SplitCLK_4_1124_DFFT_395__FPB_n1575(net1162_c1,net1162);
INTERCONNECT SplitCLK_4_1123_DFFT_459__FPB_n1639(net1163_c1,net1163);
INTERCONNECT SplitCLK_2_1122_DFFT_467__FPB_n1647(net1164_c1,net1164);
INTERCONNECT SplitCLK_2_1121_DFFT_475__FPB_n1655(net1165_c1,net1165);
INTERCONNECT SplitCLK_4_1120_DFFT_483__FPB_n1663(net1166_c1,net1166);
INTERCONNECT SplitCLK_2_1119_DFFT_491__FPB_n1671(net1167_c1,net1167);
INTERCONNECT SplitCLK_2_1118_DFFT_539__FPB_n1719(net1168_c1,net1168);
INTERCONNECT SplitCLK_4_1117_AND2T_129_n130(net1169_c1,net1169);
INTERCONNECT SplitCLK_2_1116_AND2T_118_n119(net1170_c1,net1170);
INTERCONNECT SplitCLK_2_1115_AND2T_126_n127(net1171_c1,net1171);
INTERCONNECT SplitCLK_2_1114_AND2T_141_n142(net1172_c1,net1172);
INTERCONNECT SplitCLK_2_1113_AND2T_109_n110(net1173_c1,net1173);
INTERCONNECT SplitCLK_4_1112_AND2T_116_n117(net1174_c1,net1174);
INTERCONNECT SplitCLK_4_1111_AND2T_124_n125(net1175_c1,net1175);
INTERCONNECT SplitCLK_4_1110_AND2T_132_n133(net1176_c1,net1176);
INTERCONNECT SplitCLK_4_1109_AND2T_140_n141(net1177_c1,net1177);
INTERCONNECT SplitCLK_4_1108_AND2T_123_n124(net1178_c1,net1178);
INTERCONNECT SplitCLK_4_1107_AND2T_131_n132(net1179_c1,net1179);
INTERCONNECT SplitCLK_4_1106_AND2T_106_n107(net1180_c1,net1180);
INTERCONNECT SplitCLK_4_1105_AND2T_114_n115(net1181_c1,net1181);
INTERCONNECT SplitCLK_2_1104_AND2T_112_n113(net1182_c1,net1182);
INTERCONNECT SplitCLK_2_1103_AND2T_103_n104(net1183_c1,net1183);
INTERCONNECT SplitCLK_2_1102_XOR2T_89_n90(net1184_c1,net1184);
INTERCONNECT SplitCLK_2_1101_XOR2T_93_n94(net1185_c1,net1185);
INTERCONNECT SplitCLK_4_1100_XOR2T_91_n92(net1186_c1,net1186);
INTERCONNECT SplitCLK_4_1099_XOR2T_74_n75(net1187_c1,net1187);
INTERCONNECT SplitCLK_4_1098_XOR2T_65_n66(net1188_c1,net1188);
INTERCONNECT SplitCLK_2_1097_XOR2T_72_n73(net1189_c1,net1189);
INTERCONNECT SplitCLK_2_1096_XOR2T_62_n63(net1190_c1,net1190);
INTERCONNECT SplitCLK_2_1095_XOR2T_44_n45(net1191_c1,net1191);
INTERCONNECT SplitCLK_2_1094_DFFT_298__FPB_n1478(net1192_c1,net1192);
INTERCONNECT SplitCLK_4_1093_DFFT_378__FPB_n1558(net1193_c1,net1193);
INTERCONNECT SplitCLK_2_1092_DFFT_386__FPB_n1566(net1194_c1,net1194);
INTERCONNECT SplitCLK_4_1091_DFFT_394__FPB_n1574(net1195_c1,net1195);
INTERCONNECT SplitCLK_4_1090_DFFT_458__FPB_n1638(net1196_c1,net1196);
INTERCONNECT SplitCLK_2_1089_DFFT_466__FPB_n1646(net1197_c1,net1197);
INTERCONNECT SplitCLK_4_1088_DFFT_474__FPB_n1654(net1198_c1,net1198);
INTERCONNECT SplitCLK_4_1087_DFFT_482__FPB_n1662(net1199_c1,net1199);
INTERCONNECT SplitCLK_4_1086_DFFT_490__FPB_n1670(net1200_c1,net1200);
INTERCONNECT SplitCLK_2_1085_DFFT_289__FPB_n1469(net1201_c1,net1201);
INTERCONNECT SplitCLK_4_1084_DFFT_297__FPB_n1477(net1202_c1,net1202);
INTERCONNECT SplitCLK_2_1083_DFFT_369__FPB_n1549(net1203_c1,net1203);
INTERCONNECT SplitCLK_2_1082_DFFT_377__FPB_n1557(net1204_c1,net1204);
INTERCONNECT SplitCLK_2_1081_DFFT_385__FPB_n1565(net1205_c1,net1205);
INTERCONNECT SplitCLK_2_1080_DFFT_393__FPB_n1573(net1206_c1,net1206);
INTERCONNECT SplitCLK_2_1079_DFFT_449__FPB_n1629(net1207_c1,net1207);
INTERCONNECT SplitCLK_4_1078_DFFT_457__FPB_n1637(net1208_c1,net1208);
INTERCONNECT SplitCLK_4_1077_DFFT_465__FPB_n1645(net1209_c1,net1209);
INTERCONNECT SplitCLK_4_1076_DFFT_473__FPB_n1653(net1210_c1,net1210);
INTERCONNECT SplitCLK_4_1075_DFFT_481__FPB_n1661(net1211_c1,net1211);
INTERCONNECT SplitCLK_4_1074_DFFT_529__FPB_n1709(net1212_c1,net1212);
INTERCONNECT SplitCLK_4_1073_DFFT_288__FPB_n1468(net1213_c1,net1213);
INTERCONNECT SplitCLK_4_1072_DFFT_296__FPB_n1476(net1214_c1,net1214);
INTERCONNECT SplitCLK_2_1071_DFFT_368__FPB_n1548(net1215_c1,net1215);
INTERCONNECT SplitCLK_2_1070_DFFT_376__FPB_n1556(net1216_c1,net1216);
INTERCONNECT SplitCLK_4_1069_DFFT_384__FPB_n1564(net1217_c1,net1217);
INTERCONNECT SplitCLK_4_1068_DFFT_392__FPB_n1572(net1218_c1,net1218);
INTERCONNECT SplitCLK_4_1067_DFFT_448__FPB_n1628(net1219_c1,net1219);
INTERCONNECT SplitCLK_2_1066_DFFT_456__FPB_n1636(net1220_c1,net1220);
INTERCONNECT SplitCLK_2_1065_DFFT_464__FPB_n1644(net1221_c1,net1221);
INTERCONNECT SplitCLK_4_1064_DFFT_472__FPB_n1652(net1222_c1,net1222);
INTERCONNECT SplitCLK_4_1063_DFFT_480__FPB_n1660(net1223_c1,net1223);
INTERCONNECT SplitCLK_2_1062_DFFT_528__FPB_n1708(net1224_c1,net1224);
INTERCONNECT SplitCLK_2_1061_DFFT_536__FPB_n1716(net1225_c1,net1225);
INTERCONNECT SplitCLK_4_1060_DFFT_519__FPB_n1699(net1226_c1,net1226);
INTERCONNECT SplitCLK_4_1059_DFFT_199__FPB_n1379(net1227_c1,net1227);
INTERCONNECT SplitCLK_2_1058_DFFT_279__FPB_n1459(net1228_c1,net1228);
INTERCONNECT SplitCLK_2_1057_DFFT_287__FPB_n1467(net1229_c1,net1229);
INTERCONNECT SplitCLK_4_1056_DFFT_295__FPB_n1475(net1230_c1,net1230);
INTERCONNECT SplitCLK_4_1055_DFFT_359__FPB_n1539(net1231_c1,net1231);
INTERCONNECT SplitCLK_4_1054_DFFT_367__FPB_n1547(net1232_c1,net1232);
INTERCONNECT SplitCLK_4_1053_DFFT_375__FPB_n1555(net1233_c1,net1233);
INTERCONNECT SplitCLK_2_1052_DFFT_383__FPB_n1563(net1234_c1,net1234);
INTERCONNECT SplitCLK_2_1051_DFFT_439__FPB_n1619(net1235_c1,net1235);
INTERCONNECT SplitCLK_2_1050_DFFT_447__FPB_n1627(net1236_c1,net1236);
INTERCONNECT SplitCLK_4_1049_DFFT_455__FPB_n1635(net1237_c1,net1237);
INTERCONNECT SplitCLK_4_1048_DFFT_471__FPB_n1651(net1238_c1,net1238);
INTERCONNECT SplitCLK_4_1047_DFFT_535__FPB_n1715(net1239_c1,net1239);
INTERCONNECT SplitCLK_2_1046_SplitCLK_6_915(net1240_c1,net1240);
INTERCONNECT SplitCLK_2_1046_SplitCLK_4_1045(net1241_c1,net1241);
INTERCONNECT SplitCLK_4_1045_SplitCLK_0_980(net1242_c1,net1242);
INTERCONNECT SplitCLK_4_1045_SplitCLK_2_1044(net1243_c1,net1243);
INTERCONNECT SplitCLK_2_1044_SplitCLK_6_1012(net1244_c1,net1244);
INTERCONNECT SplitCLK_2_1044_SplitCLK_4_1043(net1245_c1,net1245);
INTERCONNECT SplitCLK_4_1043_SplitCLK_0_1027(net1246_c1,net1246);
INTERCONNECT SplitCLK_4_1043_SplitCLK_2_1042(net1247_c1,net1247);
INTERCONNECT SplitCLK_2_1042_SplitCLK_6_1034(net1248_c1,net1248);
INTERCONNECT SplitCLK_2_1042_SplitCLK_4_1041(net1249_c1,net1249);
INTERCONNECT SplitCLK_4_1041_SplitCLK_4_1037(net1250_c1,net1250);
INTERCONNECT SplitCLK_4_1041_SplitCLK_2_1040(net1251_c1,net1251);
INTERCONNECT SplitCLK_2_1040_SplitCLK_6_1038(net1252_c1,net1252);
INTERCONNECT SplitCLK_2_1040_SplitCLK_4_1039(net1253_c1,net1253);
INTERCONNECT SplitCLK_4_1039_SplitCLK_2_1134(net1254_c1,net1254);
INTERCONNECT SplitCLK_4_1039_SplitCLK_4_1371(net1255_c1,net1255);
INTERCONNECT SplitCLK_6_1038_SplitCLK_4_1093(net1256_c1,net1256);
INTERCONNECT SplitCLK_6_1038_SplitCLK_2_1126(net1257_c1,net1257);
INTERCONNECT SplitCLK_4_1037_SplitCLK_4_1035(net1258_c1,net1258);
INTERCONNECT SplitCLK_4_1037_SplitCLK_4_1036(net1259_c1,net1259);
INTERCONNECT SplitCLK_4_1036_SplitCLK_2_1082(net1260_c1,net1260);
INTERCONNECT SplitCLK_4_1036_SplitCLK_4_1530(net1261_c1,net1261);
INTERCONNECT SplitCLK_4_1035_SplitCLK_4_1053(net1262_c1,net1262);
INTERCONNECT SplitCLK_4_1035_SplitCLK_2_1070(net1263_c1,net1263);
INTERCONNECT SplitCLK_6_1034_SplitCLK_0_1030(net1264_c1,net1264);
INTERCONNECT SplitCLK_6_1034_SplitCLK_6_1033(net1265_c1,net1265);
INTERCONNECT SplitCLK_6_1033_SplitCLK_6_1031(net1266_c1,net1266);
INTERCONNECT SplitCLK_6_1033_SplitCLK_4_1032(net1267_c1,net1267);
INTERCONNECT SplitCLK_4_1032_SplitCLK_4_1501(net1268_c1,net1268);
INTERCONNECT SplitCLK_4_1032_SplitCLK_2_1538(net1269_c1,net1269);
INTERCONNECT SplitCLK_6_1031_SplitCLK_2_1318(net1270_c1,net1270);
INTERCONNECT SplitCLK_6_1031_SplitCLK_4_1351(net1271_c1,net1271);
INTERCONNECT SplitCLK_0_1030_SplitCLK_6_1028(net1272_c1,net1272);
INTERCONNECT SplitCLK_0_1030_SplitCLK_4_1029(net1273_c1,net1273);
INTERCONNECT SplitCLK_4_1029_SplitCLK_4_1313(net1274_c1,net1274);
INTERCONNECT SplitCLK_4_1029_SplitCLK_2_1519(net1275_c1,net1275);
INTERCONNECT SplitCLK_6_1028_SplitCLK_2_1115(net1276_c1,net1276);
INTERCONNECT SplitCLK_6_1028_SplitCLK_4_1332(net1277_c1,net1277);
INTERCONNECT SplitCLK_0_1027_SplitCLK_6_1019(net1278_c1,net1278);
INTERCONNECT SplitCLK_0_1027_SplitCLK_4_1026(net1279_c1,net1279);
INTERCONNECT SplitCLK_4_1026_SplitCLK_0_1022(net1280_c1,net1280);
INTERCONNECT SplitCLK_4_1026_SplitCLK_2_1025(net1281_c1,net1281);
INTERCONNECT SplitCLK_2_1025_SplitCLK_0_1023(net1282_c1,net1282);
INTERCONNECT SplitCLK_2_1025_SplitCLK_6_1024(net1283_c1,net1283);
INTERCONNECT SplitCLK_6_1024_SplitCLK_4_1492(net1284_c1,net1284);
INTERCONNECT SplitCLK_6_1024_SplitCLK_2_1512(net1285_c1,net1285);
INTERCONNECT SplitCLK_0_1023_SplitCLK_4_1462(net1286_c1,net1286);
INTERCONNECT SplitCLK_0_1023_SplitCLK_2_1539(net1287_c1,net1287);
INTERCONNECT SplitCLK_0_1022_SplitCLK_6_1020(net1288_c1,net1288);
INTERCONNECT SplitCLK_0_1022_SplitCLK_4_1021(net1289_c1,net1289);
INTERCONNECT SplitCLK_4_1021_SplitCLK_4_1417(net1290_c1,net1290);
INTERCONNECT SplitCLK_4_1021_SplitCLK_2_1440(net1291_c1,net1291);
INTERCONNECT SplitCLK_6_1020_SplitCLK_4_1502(net1292_c1,net1292);
INTERCONNECT SplitCLK_6_1020_SplitCLK_2_1520(net1293_c1,net1293);
INTERCONNECT SplitCLK_6_1019_SplitCLK_4_1015(net1294_c1,net1294);
INTERCONNECT SplitCLK_6_1019_SplitCLK_2_1018(net1295_c1,net1295);
INTERCONNECT SplitCLK_2_1018_SplitCLK_6_1016(net1296_c1,net1296);
INTERCONNECT SplitCLK_2_1018_SplitCLK_4_1017(net1297_c1,net1297);
INTERCONNECT SplitCLK_4_1017_SplitCLK_2_1299(net1298_c1,net1298);
INTERCONNECT SplitCLK_4_1017_SplitCLK_4_1442(net1299_c1,net1299);
INTERCONNECT SplitCLK_6_1016_SplitCLK_4_1191(net1300_c1,net1300);
INTERCONNECT SplitCLK_6_1016_SplitCLK_2_1373(net1301_c1,net1301);
INTERCONNECT SplitCLK_4_1015_SplitCLK_0_1013(net1302_c1,net1302);
INTERCONNECT SplitCLK_4_1015_SplitCLK_2_1014(net1303_c1,net1303);
INTERCONNECT SplitCLK_2_1014_SplitCLK_2_1259(net1304_c1,net1304);
INTERCONNECT SplitCLK_2_1014_SplitCLK_4_1419(net1305_c1,net1305);
INTERCONNECT SplitCLK_0_1013_SplitCLK_4_1111(net1306_c1,net1306);
INTERCONNECT SplitCLK_0_1013_SplitCLK_2_1140(net1307_c1,net1307);
INTERCONNECT SplitCLK_6_1012_SplitCLK_0_996(net1308_c1,net1308);
INTERCONNECT SplitCLK_6_1012_SplitCLK_4_1011(net1309_c1,net1309);
INTERCONNECT SplitCLK_4_1011_SplitCLK_6_1003(net1310_c1,net1310);
INTERCONNECT SplitCLK_4_1011_SplitCLK_4_1010(net1311_c1,net1311);
INTERCONNECT SplitCLK_4_1010_SplitCLK_4_1006(net1312_c1,net1312);
INTERCONNECT SplitCLK_4_1010_SplitCLK_6_1009(net1313_c1,net1313);
INTERCONNECT SplitCLK_6_1009_SplitCLK_6_1007(net1314_c1,net1314);
INTERCONNECT SplitCLK_6_1009_SplitCLK_4_1008(net1315_c1,net1315);
INTERCONNECT SplitCLK_4_1008_SplitCLK_2_1418(net1316_c1,net1316);
INTERCONNECT SplitCLK_4_1008_SplitCLK_4_1441(net1317_c1,net1317);
INTERCONNECT SplitCLK_6_1007_SplitCLK_4_1105(net1318_c1,net1318);
INTERCONNECT SplitCLK_6_1007_SplitCLK_2_1394(net1319_c1,net1319);
INTERCONNECT SplitCLK_4_1006_SplitCLK_0_1004(net1320_c1,net1320);
INTERCONNECT SplitCLK_4_1006_SplitCLK_4_1005(net1321_c1,net1321);
INTERCONNECT SplitCLK_4_1005_SplitCLK_4_1132(net1322_c1,net1322);
INTERCONNECT SplitCLK_4_1005_SplitCLK_2_1463(net1323_c1,net1323);
INTERCONNECT SplitCLK_0_1004_SplitCLK_2_1256(net1324_c1,net1324);
INTERCONNECT SplitCLK_0_1004_SplitCLK_4_1493(net1325_c1,net1325);
INTERCONNECT SplitCLK_6_1003_SplitCLK_2_999(net1326_c1,net1326);
INTERCONNECT SplitCLK_6_1003_SplitCLK_6_1002(net1327_c1,net1327);
INTERCONNECT SplitCLK_6_1002_SplitCLK_6_1000(net1328_c1,net1328);
INTERCONNECT SplitCLK_6_1002_SplitCLK_4_1001(net1329_c1,net1329);
INTERCONNECT SplitCLK_4_1001_SplitCLK_4_1254(net1330_c1,net1330);
INTERCONNECT SplitCLK_4_1001_SplitCLK_2_1359(net1331_c1,net1331);
INTERCONNECT SplitCLK_6_1000_SplitCLK_2_1320(net1332_c1,net1332);
INTERCONNECT SplitCLK_6_1000_SplitCLK_4_1338(net1333_c1,net1333);
INTERCONNECT SplitCLK_2_999_SplitCLK_0_997(net1334_c1,net1334);
INTERCONNECT SplitCLK_2_999_SplitCLK_0_998(net1335_c1,net1335);
INTERCONNECT SplitCLK_0_998_SplitCLK_4_1054(net1336_c1,net1336);
INTERCONNECT SplitCLK_0_998_SplitCLK_2_1309(net1337_c1,net1337);
INTERCONNECT SplitCLK_0_997_SplitCLK_4_1276(net1338_c1,net1338);
INTERCONNECT SplitCLK_0_997_SplitCLK_2_1304(net1339_c1,net1339);
INTERCONNECT SplitCLK_0_996_SplitCLK_6_988(net1340_c1,net1340);
INTERCONNECT SplitCLK_0_996_SplitCLK_4_995(net1341_c1,net1341);
INTERCONNECT SplitCLK_4_995_SplitCLK_6_991(net1342_c1,net1342);
INTERCONNECT SplitCLK_4_995_SplitCLK_6_994(net1343_c1,net1343);
INTERCONNECT SplitCLK_6_994_SplitCLK_0_992(net1344_c1,net1344);
INTERCONNECT SplitCLK_6_994_SplitCLK_6_993(net1345_c1,net1345);
INTERCONNECT SplitCLK_6_993_SplitCLK_4_1108(net1346_c1,net1346);
INTERCONNECT SplitCLK_6_993_SplitCLK_4_1124(net1347_c1,net1347);
INTERCONNECT SplitCLK_0_992_SplitCLK_2_1080(net1348_c1,net1348);
INTERCONNECT SplitCLK_0_992_SplitCLK_4_1091(net1349_c1,net1349);
INTERCONNECT SplitCLK_6_991_SplitCLK_4_989(net1350_c1,net1350);
INTERCONNECT SplitCLK_6_991_SplitCLK_4_990(net1351_c1,net1351);
INTERCONNECT SplitCLK_4_990_SplitCLK_4_1145(net1352_c1,net1352);
INTERCONNECT SplitCLK_4_990_SplitCLK_4_1257(net1353_c1,net1353);
INTERCONNECT SplitCLK_4_989_SplitCLK_2_1071(net1354_c1,net1354);
INTERCONNECT SplitCLK_4_989_SplitCLK_4_1466(net1355_c1,net1355);
INTERCONNECT SplitCLK_6_988_SplitCLK_0_984(net1356_c1,net1356);
INTERCONNECT SplitCLK_6_988_SplitCLK_6_987(net1357_c1,net1357);
INTERCONNECT SplitCLK_6_987_SplitCLK_6_985(net1358_c1,net1358);
INTERCONNECT SplitCLK_6_987_SplitCLK_0_986(net1359_c1,net1359);
INTERCONNECT SplitCLK_0_986_SplitCLK_4_1266(net1360_c1,net1360);
INTERCONNECT SplitCLK_0_986_SplitCLK_4_1325(net1361_c1,net1361);
INTERCONNECT SplitCLK_6_985_SplitCLK_2_1271(net1362_c1,net1362);
INTERCONNECT SplitCLK_6_985_SplitCLK_4_1281(net1363_c1,net1363);
INTERCONNECT SplitCLK_0_984_SplitCLK_4_982(net1364_c1,net1364);
INTERCONNECT SplitCLK_0_984_SplitCLK_4_983(net1365_c1,net1365);
INTERCONNECT SplitCLK_4_983_SplitCLK_2_1097(net1366_c1,net1366);
INTERCONNECT SplitCLK_4_983_SplitCLK_2_1280(net1367_c1,net1367);
INTERCONNECT SplitCLK_4_982_SplitCLK_2_1270(net1368_c1,net1368);
INTERCONNECT SplitCLK_4_982_SplitCLK_4_981(net1369_c1,net1369);
INTERCONNECT SplitCLK_4_981_DFFT_214__FPB_n1394(net1370_c1,net1370);
INTERCONNECT SplitCLK_4_981_DFFT_231__FPB_n1411(net1371_c1,net1371);
INTERCONNECT SplitCLK_0_980_SplitCLK_6_947(net1372_c1,net1372);
INTERCONNECT SplitCLK_0_980_SplitCLK_4_979(net1373_c1,net1373);
INTERCONNECT SplitCLK_4_979_SplitCLK_0_963(net1374_c1,net1374);
INTERCONNECT SplitCLK_4_979_SplitCLK_2_978(net1375_c1,net1375);
INTERCONNECT SplitCLK_2_978_SplitCLK_6_970(net1376_c1,net1376);
INTERCONNECT SplitCLK_2_978_SplitCLK_4_977(net1377_c1,net1377);
INTERCONNECT SplitCLK_4_977_SplitCLK_4_973(net1378_c1,net1378);
INTERCONNECT SplitCLK_4_977_SplitCLK_2_976(net1379_c1,net1379);
INTERCONNECT SplitCLK_2_976_SplitCLK_6_974(net1380_c1,net1380);
INTERCONNECT SplitCLK_2_976_SplitCLK_4_975(net1381_c1,net1381);
INTERCONNECT SplitCLK_4_975_SplitCLK_4_1372(net1382_c1,net1382);
INTERCONNECT SplitCLK_4_975_SplitCLK_2_1393(net1383_c1,net1383);
INTERCONNECT SplitCLK_6_974_SplitCLK_4_1448(net1384_c1,net1384);
INTERCONNECT SplitCLK_6_974_SplitCLK_2_1478(net1385_c1,net1385);
INTERCONNECT SplitCLK_4_973_SplitCLK_4_971(net1386_c1,net1386);
INTERCONNECT SplitCLK_4_973_SplitCLK_4_972(net1387_c1,net1387);
INTERCONNECT SplitCLK_4_972_SplitCLK_2_1083(net1388_c1,net1388);
INTERCONNECT SplitCLK_4_972_SplitCLK_4_1350(net1389_c1,net1389);
INTERCONNECT SplitCLK_4_971_SplitCLK_2_1185(net1390_c1,net1390);
INTERCONNECT SplitCLK_4_971_SplitCLK_4_1189(net1391_c1,net1391);
INTERCONNECT SplitCLK_6_970_SplitCLK_6_966(net1392_c1,net1392);
INTERCONNECT SplitCLK_6_970_SplitCLK_6_969(net1393_c1,net1393);
INTERCONNECT SplitCLK_6_969_SplitCLK_6_967(net1394_c1,net1394);
INTERCONNECT SplitCLK_6_969_SplitCLK_6_968(net1395_c1,net1395);
INTERCONNECT SplitCLK_6_968_SplitCLK_4_1374(net1396_c1,net1396);
INTERCONNECT SplitCLK_6_968_SplitCLK_2_1395(net1397_c1,net1397);
INTERCONNECT SplitCLK_6_967_SplitCLK_2_1149(net1398_c1,net1398);
INTERCONNECT SplitCLK_6_967_SplitCLK_2_1464(net1399_c1,net1399);
INTERCONNECT SplitCLK_6_966_SplitCLK_4_964(net1400_c1,net1400);
INTERCONNECT SplitCLK_6_966_SplitCLK_4_965(net1401_c1,net1401);
INTERCONNECT SplitCLK_4_965_SplitCLK_4_1333(net1402_c1,net1402);
INTERCONNECT SplitCLK_4_965_SplitCLK_2_1352(net1403_c1,net1403);
INTERCONNECT SplitCLK_4_964_SplitCLK_4_1112(net1404_c1,net1404);
INTERCONNECT SplitCLK_4_964_SplitCLK_2_1260(net1405_c1,net1405);
INTERCONNECT SplitCLK_0_963_SplitCLK_6_955(net1406_c1,net1406);
INTERCONNECT SplitCLK_0_963_SplitCLK_4_962(net1407_c1,net1407);
INTERCONNECT SplitCLK_4_962_SplitCLK_0_958(net1408_c1,net1408);
INTERCONNECT SplitCLK_4_962_SplitCLK_6_961(net1409_c1,net1409);
INTERCONNECT SplitCLK_6_961_SplitCLK_6_959(net1410_c1,net1410);
INTERCONNECT SplitCLK_6_961_SplitCLK_6_960(net1411_c1,net1411);
INTERCONNECT SplitCLK_6_960_SplitCLK_4_1223(net1412_c1,net1412);
INTERCONNECT SplitCLK_6_960_SplitCLK_2_1331(net1413_c1,net1413);
INTERCONNECT SplitCLK_6_959_SplitCLK_4_1087(net1414_c1,net1414);
INTERCONNECT SplitCLK_6_959_SplitCLK_2_1300(net1415_c1,net1415);
INTERCONNECT SplitCLK_0_958_SplitCLK_6_956(net1416_c1,net1416);
INTERCONNECT SplitCLK_0_958_SplitCLK_4_957(net1417_c1,net1417);
INTERCONNECT SplitCLK_4_957_SplitCLK_2_1323(net1418_c1,net1418);
INTERCONNECT SplitCLK_4_957_SplitCLK_4_1341(net1419_c1,net1419);
INTERCONNECT SplitCLK_6_956_SplitCLK_4_1120(net1420_c1,net1420);
INTERCONNECT SplitCLK_6_956_SplitCLK_2_1284(net1421_c1,net1421);
INTERCONNECT SplitCLK_6_955_SplitCLK_4_951(net1422_c1,net1422);
INTERCONNECT SplitCLK_6_955_SplitCLK_2_954(net1423_c1,net1423);
INTERCONNECT SplitCLK_2_954_SplitCLK_0_952(net1424_c1,net1424);
INTERCONNECT SplitCLK_2_954_SplitCLK_4_953(net1425_c1,net1425);
INTERCONNECT SplitCLK_4_953_SplitCLK_2_1052(net1426_c1,net1426);
INTERCONNECT SplitCLK_4_953_SplitCLK_2_1314(net1427_c1,net1427);
INTERCONNECT SplitCLK_0_952_SplitCLK_4_1069(net1428_c1,net1428);
INTERCONNECT SplitCLK_0_952_SplitCLK_2_1252(net1429_c1,net1429);
INTERCONNECT SplitCLK_4_951_SplitCLK_0_949(net1430_c1,net1430);
INTERCONNECT SplitCLK_4_951_SplitCLK_0_950(net1431_c1,net1431);
INTERCONNECT SplitCLK_0_950_SplitCLK_2_1081(net1432_c1,net1432);
INTERCONNECT SplitCLK_0_950_SplitCLK_4_1273(net1433_c1,net1433);
INTERCONNECT SplitCLK_0_949_SplitCLK_2_1537(net1434_c1,net1434);
INTERCONNECT SplitCLK_0_949_SplitCLK_4_948(net1435_c1,net1435);
INTERCONNECT SplitCLK_4_948_DFFT_391__FPB_n1571(net1436_c1,net1436);
INTERCONNECT SplitCLK_4_948_NOTT_121_n122(net1437_c1,net1437);
INTERCONNECT SplitCLK_6_947_SplitCLK_0_931(net1438_c1,net1438);
INTERCONNECT SplitCLK_6_947_SplitCLK_2_946(net1439_c1,net1439);
INTERCONNECT SplitCLK_2_946_SplitCLK_6_938(net1440_c1,net1440);
INTERCONNECT SplitCLK_2_946_SplitCLK_4_945(net1441_c1,net1441);
INTERCONNECT SplitCLK_4_945_SplitCLK_4_941(net1442_c1,net1442);
INTERCONNECT SplitCLK_4_945_SplitCLK_6_944(net1443_c1,net1443);
INTERCONNECT SplitCLK_6_944_SplitCLK_0_942(net1444_c1,net1444);
INTERCONNECT SplitCLK_6_944_SplitCLK_6_943(net1445_c1,net1445);
INTERCONNECT SplitCLK_6_943_SplitCLK_2_1251(net1446_c1,net1446);
INTERCONNECT SplitCLK_6_943_SplitCLK_4_1508(net1447_c1,net1447);
INTERCONNECT SplitCLK_0_942_SplitCLK_4_1335(net1448_c1,net1448);
INTERCONNECT SplitCLK_0_942_SplitCLK_2_1485(net1449_c1,net1449);
INTERCONNECT SplitCLK_4_941_SplitCLK_6_939(net1450_c1,net1450);
INTERCONNECT SplitCLK_4_941_SplitCLK_4_940(net1451_c1,net1451);
INTERCONNECT SplitCLK_4_940_SplitCLK_4_1248(net1452_c1,net1452);
INTERCONNECT SplitCLK_4_940_SplitCLK_2_1354(net1453_c1,net1453);
INTERCONNECT SplitCLK_6_939_SplitCLK_4_1182(net1454_c1,net1454);
INTERCONNECT SplitCLK_6_939_SplitCLK_2_1455(net1455_c1,net1455);
INTERCONNECT SplitCLK_6_938_SplitCLK_4_934(net1456_c1,net1456);
INTERCONNECT SplitCLK_6_938_SplitCLK_2_937(net1457_c1,net1457);
INTERCONNECT SplitCLK_2_937_SplitCLK_6_935(net1458_c1,net1458);
INTERCONNECT SplitCLK_2_937_SplitCLK_4_936(net1459_c1,net1459);
INTERCONNECT SplitCLK_4_936_SplitCLK_4_1208(net1460_c1,net1460);
INTERCONNECT SplitCLK_4_936_SplitCLK_2_1287(net1461_c1,net1461);
INTERCONNECT SplitCLK_6_935_SplitCLK_2_1230(net1462_c1,net1462);
INTERCONNECT SplitCLK_6_935_SplitCLK_4_1316(net1463_c1,net1463);
INTERCONNECT SplitCLK_4_934_SplitCLK_0_932(net1464_c1,net1464);
INTERCONNECT SplitCLK_4_934_SplitCLK_2_933(net1465_c1,net1465);
INTERCONNECT SplitCLK_2_933_SplitCLK_2_1243(net1466_c1,net1466);
INTERCONNECT SplitCLK_2_933_SplitCLK_4_1289(net1467_c1,net1467);
INTERCONNECT SplitCLK_0_932_SplitCLK_2_1286(net1468_c1,net1468);
INTERCONNECT SplitCLK_0_932_SplitCLK_4_1522(net1469_c1,net1469);
INTERCONNECT SplitCLK_0_931_SplitCLK_6_923(net1470_c1,net1470);
INTERCONNECT SplitCLK_0_931_SplitCLK_4_930(net1471_c1,net1471);
INTERCONNECT SplitCLK_4_930_SplitCLK_0_926(net1472_c1,net1472);
INTERCONNECT SplitCLK_4_930_SplitCLK_6_929(net1473_c1,net1473);
INTERCONNECT SplitCLK_6_929_SplitCLK_0_927(net1474_c1,net1474);
INTERCONNECT SplitCLK_6_929_SplitCLK_6_928(net1475_c1,net1475);
INTERCONNECT SplitCLK_6_928_SplitCLK_4_1178(net1476_c1,net1476);
INTERCONNECT SplitCLK_6_928_SplitCLK_2_1179(net1477_c1,net1477);
INTERCONNECT SplitCLK_0_927_SplitCLK_2_1116(net1478_c1,net1478);
INTERCONNECT SplitCLK_0_927_SplitCLK_4_1125(net1479_c1,net1479);
INTERCONNECT SplitCLK_0_926_SplitCLK_6_924(net1480_c1,net1480);
INTERCONNECT SplitCLK_0_926_SplitCLK_0_925(net1481_c1,net1481);
INTERCONNECT SplitCLK_0_925_SplitCLK_2_1133(net1482_c1,net1482);
INTERCONNECT SplitCLK_0_925_SplitCLK_4_1210(net1483_c1,net1483);
INTERCONNECT SplitCLK_6_924_SplitCLK_2_1521(net1484_c1,net1484);
INTERCONNECT SplitCLK_6_924_SplitCLK_4_1540(net1485_c1,net1485);
INTERCONNECT SplitCLK_6_923_SplitCLK_6_919(net1486_c1,net1486);
INTERCONNECT SplitCLK_6_923_SplitCLK_2_922(net1487_c1,net1487);
INTERCONNECT SplitCLK_2_922_SplitCLK_6_920(net1488_c1,net1488);
INTERCONNECT SplitCLK_2_922_SplitCLK_4_921(net1489_c1,net1489);
INTERCONNECT SplitCLK_4_921_SplitCLK_2_1092(net1490_c1,net1490);
INTERCONNECT SplitCLK_4_921_SplitCLK_2_1218(net1491_c1,net1491);
INTERCONNECT SplitCLK_6_920_SplitCLK_2_1113(net1492_c1,net1492);
INTERCONNECT SplitCLK_6_920_SplitCLK_2_1404(net1493_c1,net1493);
INTERCONNECT SplitCLK_6_919_SplitCLK_4_917(net1494_c1,net1494);
INTERCONNECT SplitCLK_6_919_SplitCLK_4_918(net1495_c1,net1495);
INTERCONNECT SplitCLK_4_918_SplitCLK_4_1233(net1496_c1,net1496);
INTERCONNECT SplitCLK_4_918_SplitCLK_2_1253(net1497_c1,net1497);
INTERCONNECT SplitCLK_4_917_SplitCLK_2_1258(net1498_c1,net1498);
INTERCONNECT SplitCLK_4_917_SplitCLK_4_916(net1499_c1,net1499);
INTERCONNECT SplitCLK_4_916_OR2T_111_n112(net1500_c1,net1500);
INTERCONNECT SplitCLK_4_916_DFFT_353__FPB_n1533(net1501_c1,net1501);
INTERCONNECT SplitCLK_6_915_SplitCLK_6_850(net1502_c1,net1502);
INTERCONNECT SplitCLK_6_915_SplitCLK_2_914(net1503_c1,net1503);
INTERCONNECT SplitCLK_2_914_SplitCLK_6_882(net1504_c1,net1504);
INTERCONNECT SplitCLK_2_914_SplitCLK_4_913(net1505_c1,net1505);
INTERCONNECT SplitCLK_4_913_SplitCLK_0_897(net1506_c1,net1506);
INTERCONNECT SplitCLK_4_913_SplitCLK_2_912(net1507_c1,net1507);
INTERCONNECT SplitCLK_2_912_SplitCLK_6_904(net1508_c1,net1508);
INTERCONNECT SplitCLK_2_912_SplitCLK_4_911(net1509_c1,net1509);
INTERCONNECT SplitCLK_4_911_SplitCLK_4_907(net1510_c1,net1510);
INTERCONNECT SplitCLK_4_911_SplitCLK_2_910(net1511_c1,net1511);
INTERCONNECT SplitCLK_2_910_SplitCLK_6_908(net1512_c1,net1512);
INTERCONNECT SplitCLK_2_910_SplitCLK_4_909(net1513_c1,net1513);
INTERCONNECT SplitCLK_4_909_SplitCLK_4_1290(net1514_c1,net1514);
INTERCONNECT SplitCLK_4_909_SplitCLK_2_1429(net1515_c1,net1515);
INTERCONNECT SplitCLK_6_908_SplitCLK_2_1360(net1516_c1,net1516);
INTERCONNECT SplitCLK_6_908_SplitCLK_4_1407(net1517_c1,net1517);
INTERCONNECT SplitCLK_4_907_SplitCLK_0_905(net1518_c1,net1518);
INTERCONNECT SplitCLK_4_907_SplitCLK_4_906(net1519_c1,net1519);
INTERCONNECT SplitCLK_4_906_SplitCLK_4_1228(net1520_c1,net1520);
INTERCONNECT SplitCLK_4_906_SplitCLK_2_1382(net1521_c1,net1521);
INTERCONNECT SplitCLK_0_905_SplitCLK_4_1246(net1522_c1,net1522);
INTERCONNECT SplitCLK_0_905_SplitCLK_2_1339(net1523_c1,net1523);
INTERCONNECT SplitCLK_6_904_SplitCLK_0_900(net1524_c1,net1524);
INTERCONNECT SplitCLK_6_904_SplitCLK_6_903(net1525_c1,net1525);
INTERCONNECT SplitCLK_6_903_SplitCLK_6_901(net1526_c1,net1526);
INTERCONNECT SplitCLK_6_903_SplitCLK_4_902(net1527_c1,net1527);
INTERCONNECT SplitCLK_4_902_SplitCLK_2_1236(net1528_c1,net1528);
INTERCONNECT SplitCLK_4_902_SplitCLK_4_1303(net1529_c1,net1529);
INTERCONNECT SplitCLK_6_901_SplitCLK_2_1058(net1530_c1,net1530);
INTERCONNECT SplitCLK_6_901_SplitCLK_4_1544(net1531_c1,net1531);
INTERCONNECT SplitCLK_0_900_SplitCLK_0_898(net1532_c1,net1532);
INTERCONNECT SplitCLK_0_900_SplitCLK_4_899(net1533_c1,net1533);
INTERCONNECT SplitCLK_4_899_SplitCLK_4_1224(net1534_c1,net1534);
INTERCONNECT SplitCLK_4_899_SplitCLK_2_1317(net1535_c1,net1535);
INTERCONNECT SplitCLK_0_898_SplitCLK_4_1075(net1536_c1,net1536);
INTERCONNECT SplitCLK_0_898_SplitCLK_2_1102(net1537_c1,net1537);
INTERCONNECT SplitCLK_0_897_SplitCLK_6_889(net1538_c1,net1538);
INTERCONNECT SplitCLK_0_897_SplitCLK_4_896(net1539_c1,net1539);
INTERCONNECT SplitCLK_4_896_SplitCLK_0_892(net1540_c1,net1540);
INTERCONNECT SplitCLK_4_896_SplitCLK_6_895(net1541_c1,net1541);
INTERCONNECT SplitCLK_6_895_SplitCLK_2_893(net1542_c1,net1542);
INTERCONNECT SplitCLK_6_895_SplitCLK_4_894(net1543_c1,net1543);
INTERCONNECT SplitCLK_4_894_SplitCLK_2_1263(net1544_c1,net1544);
INTERCONNECT SplitCLK_4_894_SplitCLK_4_1295(net1545_c1,net1545);
INTERCONNECT SplitCLK_2_893_SplitCLK_4_1187(net1546_c1,net1546);
INTERCONNECT SplitCLK_2_893_SplitCLK_2_1277(net1547_c1,net1547);
INTERCONNECT SplitCLK_0_892_SplitCLK_6_890(net1548_c1,net1548);
INTERCONNECT SplitCLK_0_892_SplitCLK_0_891(net1549_c1,net1549);
INTERCONNECT SplitCLK_0_891_SplitCLK_2_1221(net1550_c1,net1550);
INTERCONNECT SplitCLK_0_891_SplitCLK_4_1226(net1551_c1,net1551);
INTERCONNECT SplitCLK_6_890_SplitCLK_4_1225(net1552_c1,net1552);
INTERCONNECT SplitCLK_6_890_SplitCLK_2_1288(net1553_c1,net1553);
INTERCONNECT SplitCLK_6_889_SplitCLK_4_885(net1554_c1,net1554);
INTERCONNECT SplitCLK_6_889_SplitCLK_2_888(net1555_c1,net1555);
INTERCONNECT SplitCLK_2_888_SplitCLK_6_886(net1556_c1,net1556);
INTERCONNECT SplitCLK_2_888_SplitCLK_4_887(net1557_c1,net1557);
INTERCONNECT SplitCLK_4_887_SplitCLK_4_1063(net1558_c1,net1558);
INTERCONNECT SplitCLK_4_887_SplitCLK_2_1267(net1559_c1,net1559);
INTERCONNECT SplitCLK_6_886_SplitCLK_4_1397(net1560_c1,net1560);
INTERCONNECT SplitCLK_6_886_SplitCLK_2_1454(net1561_c1,net1561);
INTERCONNECT SplitCLK_4_885_SplitCLK_0_883(net1562_c1,net1562);
INTERCONNECT SplitCLK_4_885_SplitCLK_4_884(net1563_c1,net1563);
INTERCONNECT SplitCLK_4_884_SplitCLK_4_1144(net1564_c1,net1564);
INTERCONNECT SplitCLK_4_884_SplitCLK_2_1148(net1565_c1,net1565);
INTERCONNECT SplitCLK_0_883_SplitCLK_4_1415(net1566_c1,net1566);
INTERCONNECT SplitCLK_0_883_SplitCLK_2_1438(net1567_c1,net1567);
INTERCONNECT SplitCLK_6_882_SplitCLK_0_866(net1568_c1,net1568);
INTERCONNECT SplitCLK_6_882_SplitCLK_2_881(net1569_c1,net1569);
INTERCONNECT SplitCLK_2_881_SplitCLK_6_873(net1570_c1,net1570);
INTERCONNECT SplitCLK_2_881_SplitCLK_4_880(net1571_c1,net1571);
INTERCONNECT SplitCLK_4_880_SplitCLK_4_876(net1572_c1,net1572);
INTERCONNECT SplitCLK_4_880_SplitCLK_2_879(net1573_c1,net1573);
INTERCONNECT SplitCLK_2_879_SplitCLK_0_877(net1574_c1,net1574);
INTERCONNECT SplitCLK_2_879_SplitCLK_0_878(net1575_c1,net1575);
INTERCONNECT SplitCLK_0_878_SplitCLK_4_1408(net1576_c1,net1576);
INTERCONNECT SplitCLK_0_878_SplitCLK_2_1507(net1577_c1,net1577);
INTERCONNECT SplitCLK_0_877_SplitCLK_2_1272(net1578_c1,net1578);
INTERCONNECT SplitCLK_0_877_SplitCLK_4_1282(net1579_c1,net1579);
INTERCONNECT SplitCLK_4_876_SplitCLK_6_874(net1580_c1,net1580);
INTERCONNECT SplitCLK_4_876_SplitCLK_0_875(net1581_c1,net1581);
INTERCONNECT SplitCLK_0_875_SplitCLK_2_1215(net1582_c1,net1582);
INTERCONNECT SplitCLK_0_875_SplitCLK_4_1430(net1583_c1,net1583);
INTERCONNECT SplitCLK_6_874_SplitCLK_4_1330(net1584_c1,net1584);
INTERCONNECT SplitCLK_6_874_SplitCLK_2_1398(net1585_c1,net1585);
INTERCONNECT SplitCLK_6_873_SplitCLK_0_869(net1586_c1,net1586);
INTERCONNECT SplitCLK_6_873_SplitCLK_6_872(net1587_c1,net1587);
INTERCONNECT SplitCLK_6_872_SplitCLK_6_870(net1588_c1,net1588);
INTERCONNECT SplitCLK_6_872_SplitCLK_4_871(net1589_c1,net1589);
INTERCONNECT SplitCLK_4_871_SplitCLK_4_1392(net1590_c1,net1590);
INTERCONNECT SplitCLK_4_871_SplitCLK_2_1511(net1591_c1,net1591);
INTERCONNECT SplitCLK_6_870_SplitCLK_4_1491(net1592_c1,net1592);
INTERCONNECT SplitCLK_6_870_SplitCLK_2_1529(net1593_c1,net1593);
INTERCONNECT SplitCLK_0_869_SplitCLK_6_867(net1594_c1,net1594);
INTERCONNECT SplitCLK_0_869_SplitCLK_0_868(net1595_c1,net1595);
INTERCONNECT SplitCLK_0_868_SplitCLK_4_1370(net1596_c1,net1596);
INTERCONNECT SplitCLK_0_868_SplitCLK_2_1461(net1597_c1,net1597);
INTERCONNECT SplitCLK_6_867_SplitCLK_4_1060(net1598_c1,net1598);
INTERCONNECT SplitCLK_6_867_SplitCLK_2_1546(net1599_c1,net1599);
INTERCONNECT SplitCLK_0_866_SplitCLK_6_858(net1600_c1,net1600);
INTERCONNECT SplitCLK_0_866_SplitCLK_4_865(net1601_c1,net1601);
INTERCONNECT SplitCLK_4_865_SplitCLK_4_861(net1602_c1,net1602);
INTERCONNECT SplitCLK_4_865_SplitCLK_6_864(net1603_c1,net1603);
INTERCONNECT SplitCLK_6_864_SplitCLK_4_862(net1604_c1,net1604);
INTERCONNECT SplitCLK_6_864_SplitCLK_6_863(net1605_c1,net1605);
INTERCONNECT SplitCLK_6_863_SplitCLK_4_1327(net1606_c1,net1606);
INTERCONNECT SplitCLK_6_863_SplitCLK_2_1484(net1607_c1,net1607);
INTERCONNECT SplitCLK_4_862_SplitCLK_2_1156(net1608_c1,net1608);
INTERCONNECT SplitCLK_4_862_SplitCLK_2_1346(net1609_c1,net1609);
INTERCONNECT SplitCLK_4_861_SplitCLK_6_859(net1610_c1,net1610);
INTERCONNECT SplitCLK_4_861_SplitCLK_4_860(net1611_c1,net1611);
INTERCONNECT SplitCLK_4_860_SplitCLK_4_1296(net1612_c1,net1612);
INTERCONNECT SplitCLK_4_860_SplitCLK_2_1368(net1613_c1,net1613);
INTERCONNECT SplitCLK_6_859_SplitCLK_4_1155(net1614_c1,net1614);
INTERCONNECT SplitCLK_6_859_SplitCLK_4_1204(net1615_c1,net1615);
INTERCONNECT SplitCLK_6_858_SplitCLK_6_854(net1616_c1,net1616);
INTERCONNECT SplitCLK_6_858_SplitCLK_2_857(net1617_c1,net1617);
INTERCONNECT SplitCLK_2_857_SplitCLK_6_855(net1618_c1,net1618);
INTERCONNECT SplitCLK_2_857_SplitCLK_0_856(net1619_c1,net1619);
INTERCONNECT SplitCLK_0_856_SplitCLK_4_1198(net1620_c1,net1620);
INTERCONNECT SplitCLK_0_856_SplitCLK_2_1469(net1621_c1,net1621);
INTERCONNECT SplitCLK_6_855_SplitCLK_2_1399(net1622_c1,net1622);
INTERCONNECT SplitCLK_6_855_SplitCLK_4_1439(net1623_c1,net1623);
INTERCONNECT SplitCLK_6_854_SplitCLK_4_852(net1624_c1,net1624);
INTERCONNECT SplitCLK_6_854_SplitCLK_4_853(net1625_c1,net1625);
INTERCONNECT SplitCLK_4_853_SplitCLK_4_1160(net1626_c1,net1626);
INTERCONNECT SplitCLK_4_853_SplitCLK_2_1416(net1627_c1,net1627);
INTERCONNECT SplitCLK_4_852_SplitCLK_2_1422(net1628_c1,net1628);
INTERCONNECT SplitCLK_4_852_SplitCLK_4_851(net1629_c1,net1629);
INTERCONNECT SplitCLK_4_851_DFFT_537__FPB_n1717(net1630_c1,net1630);
INTERCONNECT SplitCLK_4_851_DFFT_522__FPB_n1702(net1631_c1,net1631);
INTERCONNECT SplitCLK_6_850_SplitCLK_6_817(net1632_c1,net1632);
INTERCONNECT SplitCLK_6_850_SplitCLK_4_849(net1633_c1,net1633);
INTERCONNECT SplitCLK_4_849_SplitCLK_0_833(net1634_c1,net1634);
INTERCONNECT SplitCLK_4_849_SplitCLK_4_848(net1635_c1,net1635);
INTERCONNECT SplitCLK_4_848_SplitCLK_6_840(net1636_c1,net1636);
INTERCONNECT SplitCLK_4_848_SplitCLK_4_847(net1637_c1,net1637);
INTERCONNECT SplitCLK_4_847_SplitCLK_0_843(net1638_c1,net1638);
INTERCONNECT SplitCLK_4_847_SplitCLK_6_846(net1639_c1,net1639);
INTERCONNECT SplitCLK_6_846_SplitCLK_6_844(net1640_c1,net1640);
INTERCONNECT SplitCLK_6_846_SplitCLK_4_845(net1641_c1,net1641);
INTERCONNECT SplitCLK_4_845_SplitCLK_2_1249(net1642_c1,net1642);
INTERCONNECT SplitCLK_4_845_SplitCLK_4_1265(net1643_c1,net1643);
INTERCONNECT SplitCLK_6_844_SplitCLK_4_1072(net1644_c1,net1644);
INTERCONNECT SplitCLK_6_844_SplitCLK_2_1229(net1645_c1,net1645);
INTERCONNECT SplitCLK_0_843_SplitCLK_6_841(net1646_c1,net1646);
INTERCONNECT SplitCLK_0_843_SplitCLK_4_842(net1647_c1,net1647);
INTERCONNECT SplitCLK_4_842_SplitCLK_2_1275(net1648_c1,net1648);
INTERCONNECT SplitCLK_4_842_SplitCLK_4_1302(net1649_c1,net1649);
INTERCONNECT SplitCLK_6_841_SplitCLK_2_1094(net1650_c1,net1650);
INTERCONNECT SplitCLK_6_841_SplitCLK_4_1220(net1651_c1,net1651);
INTERCONNECT SplitCLK_6_840_SplitCLK_0_836(net1652_c1,net1652);
INTERCONNECT SplitCLK_6_840_SplitCLK_6_839(net1653_c1,net1653);
INTERCONNECT SplitCLK_6_839_SplitCLK_2_837(net1654_c1,net1654);
INTERCONNECT SplitCLK_6_839_SplitCLK_4_838(net1655_c1,net1655);
INTERCONNECT SplitCLK_4_838_SplitCLK_4_1084(net1656_c1,net1656);
INTERCONNECT SplitCLK_4_838_SplitCLK_2_1127(net1657_c1,net1657);
INTERCONNECT SplitCLK_2_837_SplitCLK_4_1139(net1658_c1,net1658);
INTERCONNECT SplitCLK_2_837_SplitCLK_2_1468(net1659_c1,net1659);
INTERCONNECT SplitCLK_0_836_SplitCLK_6_834(net1660_c1,net1660);
INTERCONNECT SplitCLK_0_836_SplitCLK_4_835(net1661_c1,net1661);
INTERCONNECT SplitCLK_4_835_SplitCLK_2_1244(net1662_c1,net1662);
INTERCONNECT SplitCLK_4_835_SplitCLK_4_1451(net1663_c1,net1663);
INTERCONNECT SplitCLK_6_834_SplitCLK_4_1056(net1664_c1,net1664);
INTERCONNECT SplitCLK_6_834_SplitCLK_2_1219(net1665_c1,net1665);
INTERCONNECT SplitCLK_0_833_SplitCLK_4_825(net1666_c1,net1666);
INTERCONNECT SplitCLK_0_833_SplitCLK_4_832(net1667_c1,net1667);
INTERCONNECT SplitCLK_4_832_SplitCLK_0_828(net1668_c1,net1668);
INTERCONNECT SplitCLK_4_832_SplitCLK_2_831(net1669_c1,net1669);
INTERCONNECT SplitCLK_2_831_SplitCLK_6_829(net1670_c1,net1670);
INTERCONNECT SplitCLK_2_831_SplitCLK_4_830(net1671_c1,net1671);
INTERCONNECT SplitCLK_4_830_SplitCLK_2_1173(net1672_c1,net1672);
INTERCONNECT SplitCLK_4_830_SplitCLK_4_1379(net1673_c1,net1673);
INTERCONNECT SplitCLK_6_829_SplitCLK_2_1345(net1674_c1,net1674);
INTERCONNECT SplitCLK_6_829_SplitCLK_4_1367(net1675_c1,net1675);
INTERCONNECT SplitCLK_0_828_SplitCLK_4_826(net1676_c1,net1676);
INTERCONNECT SplitCLK_0_828_SplitCLK_4_827(net1677_c1,net1677);
INTERCONNECT SplitCLK_4_827_SplitCLK_2_1481(net1678_c1,net1678);
INTERCONNECT SplitCLK_4_827_SplitCLK_4_1505(net1679_c1,net1679);
INTERCONNECT SplitCLK_4_826_SplitCLK_2_1389(net1680_c1,net1680);
INTERCONNECT SplitCLK_4_826_SplitCLK_4_1413(net1681_c1,net1681);
INTERCONNECT SplitCLK_4_825_SplitCLK_0_821(net1682_c1,net1682);
INTERCONNECT SplitCLK_4_825_SplitCLK_6_824(net1683_c1,net1683);
INTERCONNECT SplitCLK_6_824_SplitCLK_4_822(net1684_c1,net1684);
INTERCONNECT SplitCLK_6_824_SplitCLK_4_823(net1685_c1,net1685);
INTERCONNECT SplitCLK_4_823_SplitCLK_4_1109(net1686_c1,net1686);
INTERCONNECT SplitCLK_4_823_SplitCLK_2_1161(net1687_c1,net1687);
INTERCONNECT SplitCLK_4_822_SplitCLK_2_1101(net1688_c1,net1688);
INTERCONNECT SplitCLK_4_822_SplitCLK_2_1157(net1689_c1,net1689);
INTERCONNECT SplitCLK_0_821_SplitCLK_2_819(net1690_c1,net1690);
INTERCONNECT SplitCLK_0_821_SplitCLK_4_820(net1691_c1,net1691);
INTERCONNECT SplitCLK_4_820_SplitCLK_4_1175(net1692_c1,net1692);
INTERCONNECT SplitCLK_4_820_SplitCLK_2_1193(net1693_c1,net1693);
INTERCONNECT SplitCLK_2_819_SplitCLK_2_1194(net1694_c1,net1694);
INTERCONNECT SplitCLK_2_819_SplitCLK_4_818(net1695_c1,net1695);
INTERCONNECT SplitCLK_4_818_DFFT_151__FPB_n1331(net1696_c1,net1696);
INTERCONNECT SplitCLK_4_818_DFFT_152__FPB_n1332(net1697_c1,net1697);
INTERCONNECT SplitCLK_6_817_SplitCLK_0_801(net1698_c1,net1698);
INTERCONNECT SplitCLK_6_817_SplitCLK_2_816(net1699_c1,net1699);
INTERCONNECT SplitCLK_2_816_SplitCLK_6_808(net1700_c1,net1700);
INTERCONNECT SplitCLK_2_816_SplitCLK_4_815(net1701_c1,net1701);
INTERCONNECT SplitCLK_4_815_SplitCLK_4_811(net1702_c1,net1702);
INTERCONNECT SplitCLK_4_815_SplitCLK_2_814(net1703_c1,net1703);
INTERCONNECT SplitCLK_2_814_SplitCLK_6_812(net1704_c1,net1704);
INTERCONNECT SplitCLK_2_814_SplitCLK_4_813(net1705_c1,net1705);
INTERCONNECT SplitCLK_4_813_SplitCLK_2_1095(net1706_c1,net1706);
INTERCONNECT SplitCLK_4_813_SplitCLK_2_1310(net1707_c1,net1707);
INTERCONNECT SplitCLK_6_812_SplitCLK_2_1158(net1708_c1,net1708);
INTERCONNECT SplitCLK_6_812_SplitCLK_2_1391(net1709_c1,net1709);
INTERCONNECT SplitCLK_4_811_SplitCLK_6_809(net1710_c1,net1710);
INTERCONNECT SplitCLK_4_811_SplitCLK_4_810(net1711_c1,net1711);
INTERCONNECT SplitCLK_4_810_SplitCLK_2_1152(net1712_c1,net1712);
INTERCONNECT SplitCLK_4_810_SplitCLK_4_1349(net1713_c1,net1713);
INTERCONNECT SplitCLK_6_809_SplitCLK_4_1100(net1714_c1,net1714);
INTERCONNECT SplitCLK_6_809_SplitCLK_2_1151(net1715_c1,net1715);
INTERCONNECT SplitCLK_6_808_SplitCLK_0_804(net1716_c1,net1716);
INTERCONNECT SplitCLK_6_808_SplitCLK_6_807(net1717_c1,net1717);
INTERCONNECT SplitCLK_6_807_SplitCLK_6_805(net1718_c1,net1718);
INTERCONNECT SplitCLK_6_807_SplitCLK_6_806(net1719_c1,net1719);
INTERCONNECT SplitCLK_6_806_SplitCLK_4_1206(net1720_c1,net1720);
INTERCONNECT SplitCLK_6_806_SplitCLK_2_1247(net1721_c1,net1721);
INTERCONNECT SplitCLK_6_805_SplitCLK_4_1047(net1722_c1,net1722);
INTERCONNECT SplitCLK_6_805_SplitCLK_2_1061(net1723_c1,net1723);
INTERCONNECT SplitCLK_0_804_SplitCLK_6_802(net1724_c1,net1724);
INTERCONNECT SplitCLK_0_804_SplitCLK_0_803(net1725_c1,net1725);
INTERCONNECT SplitCLK_0_803_SplitCLK_4_1195(net1726_c1,net1726);
INTERCONNECT SplitCLK_0_803_SplitCLK_2_1437(net1727_c1,net1727);
INTERCONNECT SplitCLK_6_802_SplitCLK_4_1513(net1728_c1,net1728);
INTERCONNECT SplitCLK_6_802_SplitCLK_2_1531(net1729_c1,net1729);
INTERCONNECT SplitCLK_0_801_SplitCLK_6_793(net1730_c1,net1730);
INTERCONNECT SplitCLK_0_801_SplitCLK_4_800(net1731_c1,net1731);
INTERCONNECT SplitCLK_4_800_SplitCLK_0_796(net1732_c1,net1732);
INTERCONNECT SplitCLK_4_800_SplitCLK_2_799(net1733_c1,net1733);
INTERCONNECT SplitCLK_2_799_SplitCLK_6_797(net1734_c1,net1734);
INTERCONNECT SplitCLK_2_799_SplitCLK_4_798(net1735_c1,net1735);
INTERCONNECT SplitCLK_4_798_SplitCLK_2_1180(net1736_c1,net1736);
INTERCONNECT SplitCLK_4_798_SplitCLK_4_1525(net1737_c1,net1737);
INTERCONNECT SplitCLK_6_797_SplitCLK_4_1192(net1738_c1,net1738);
INTERCONNECT SplitCLK_6_797_SplitCLK_2_1196(net1739_c1,net1739);
INTERCONNECT SplitCLK_0_796_SplitCLK_4_794(net1740_c1,net1740);
INTERCONNECT SplitCLK_0_796_SplitCLK_4_795(net1741_c1,net1741);
INTERCONNECT SplitCLK_4_795_SplitCLK_4_1200(net1742_c1,net1742);
INTERCONNECT SplitCLK_4_795_SplitCLK_2_1526(net1743_c1,net1743);
INTERCONNECT SplitCLK_4_794_SplitCLK_2_1197(net1744_c1,net1744);
INTERCONNECT SplitCLK_4_794_SplitCLK_2_1458(net1745_c1,net1745);
INTERCONNECT SplitCLK_6_793_SplitCLK_4_789(net1746_c1,net1746);
INTERCONNECT SplitCLK_6_793_SplitCLK_6_792(net1747_c1,net1747);
INTERCONNECT SplitCLK_6_792_SplitCLK_6_790(net1748_c1,net1748);
INTERCONNECT SplitCLK_6_792_SplitCLK_6_791(net1749_c1,net1749);
INTERCONNECT SplitCLK_6_791_SplitCLK_4_1390(net1750_c1,net1750);
INTERCONNECT SplitCLK_6_791_SplitCLK_2_1414(net1751_c1,net1751);
INTERCONNECT SplitCLK_6_790_SplitCLK_4_1472(net1752_c1,net1752);
INTERCONNECT SplitCLK_6_790_SplitCLK_2_1494(net1753_c1,net1753);
INTERCONNECT SplitCLK_4_789_SplitCLK_2_787(net1754_c1,net1754);
INTERCONNECT SplitCLK_4_789_SplitCLK_2_788(net1755_c1,net1755);
INTERCONNECT SplitCLK_2_788_SplitCLK_2_1162(net1756_c1,net1756);
INTERCONNECT SplitCLK_2_788_SplitCLK_4_1435(net1757_c1,net1757);
INTERCONNECT SplitCLK_2_787_SplitCLK_2_1135(net1758_c1,net1758);
INTERCONNECT SplitCLK_2_787_SplitCLK_4_786(net1759_c1,net1759);
INTERCONNECT SplitCLK_4_786_DFFT_538_Q1(net1760_c1,net1760);
INTERCONNECT SplitCLK_4_786_DFFT_192__FPB_n1372(net1761_c1,net1761);
INTERCONNECT SplitCLK_0_785_SplitCLK_6_654(net1762_c1,net1762);
INTERCONNECT SplitCLK_0_785_SplitCLK_4_784(net1763_c1,net1763);
INTERCONNECT SplitCLK_4_784_SplitCLK_0_719(net1764_c1,net1764);
INTERCONNECT SplitCLK_4_784_SplitCLK_4_783(net1765_c1,net1765);
INTERCONNECT SplitCLK_4_783_SplitCLK_6_751(net1766_c1,net1766);
INTERCONNECT SplitCLK_4_783_SplitCLK_4_782(net1767_c1,net1767);
INTERCONNECT SplitCLK_4_782_SplitCLK_0_766(net1768_c1,net1768);
INTERCONNECT SplitCLK_4_782_SplitCLK_6_781(net1769_c1,net1769);
INTERCONNECT SplitCLK_6_781_SplitCLK_4_773(net1770_c1,net1770);
INTERCONNECT SplitCLK_6_781_SplitCLK_4_780(net1771_c1,net1771);
INTERCONNECT SplitCLK_4_780_SplitCLK_0_776(net1772_c1,net1772);
INTERCONNECT SplitCLK_4_780_SplitCLK_2_779(net1773_c1,net1773);
INTERCONNECT SplitCLK_2_779_SplitCLK_6_777(net1774_c1,net1774);
INTERCONNECT SplitCLK_2_779_SplitCLK_4_778(net1775_c1,net1775);
INTERCONNECT SplitCLK_4_778_SplitCLK_2_1423(net1776_c1,net1776);
INTERCONNECT SplitCLK_4_778_SplitCLK_4_1445(net1777_c1,net1777);
INTERCONNECT SplitCLK_6_777_SplitCLK_2_1129(net1778_c1,net1778);
INTERCONNECT SplitCLK_6_777_SplitCLK_4_1138(net1779_c1,net1779);
INTERCONNECT SplitCLK_0_776_SplitCLK_4_774(net1780_c1,net1780);
INTERCONNECT SplitCLK_0_776_SplitCLK_4_775(net1781_c1,net1781);
INTERCONNECT SplitCLK_4_775_SplitCLK_2_1475(net1782_c1,net1782);
INTERCONNECT SplitCLK_4_775_SplitCLK_4_1498(net1783_c1,net1783);
INTERCONNECT SplitCLK_4_774_SplitCLK_2_1143(net1784_c1,net1784);
INTERCONNECT SplitCLK_4_774_SplitCLK_4_1147(net1785_c1,net1785);
INTERCONNECT SplitCLK_4_773_SplitCLK_6_769(net1786_c1,net1786);
INTERCONNECT SplitCLK_4_773_SplitCLK_6_772(net1787_c1,net1787);
INTERCONNECT SplitCLK_6_772_SplitCLK_6_770(net1788_c1,net1788);
INTERCONNECT SplitCLK_6_772_SplitCLK_6_771(net1789_c1,net1789);
INTERCONNECT SplitCLK_6_771_SplitCLK_2_1238(net1790_c1,net1790);
INTERCONNECT SplitCLK_6_771_SplitCLK_4_1543(net1791_c1,net1791);
INTERCONNECT SplitCLK_6_770_SplitCLK_4_1068(net1792_c1,net1792);
INTERCONNECT SplitCLK_6_770_SplitCLK_2_1150(net1793_c1,net1793);
INTERCONNECT SplitCLK_6_769_SplitCLK_4_767(net1794_c1,net1794);
INTERCONNECT SplitCLK_6_769_SplitCLK_4_768(net1795_c1,net1795);
INTERCONNECT SplitCLK_4_768_SplitCLK_2_1057(net1796_c1,net1796);
INTERCONNECT SplitCLK_4_768_SplitCLK_4_1073(net1797_c1,net1797);
INTERCONNECT SplitCLK_4_767_SplitCLK_2_1261(net1798_c1,net1798);
INTERCONNECT SplitCLK_4_767_SplitCLK_4_1524(net1799_c1,net1799);
INTERCONNECT SplitCLK_0_766_SplitCLK_6_758(net1800_c1,net1800);
INTERCONNECT SplitCLK_0_766_SplitCLK_4_765(net1801_c1,net1801);
INTERCONNECT SplitCLK_4_765_SplitCLK_0_761(net1802_c1,net1802);
INTERCONNECT SplitCLK_4_765_SplitCLK_4_764(net1803_c1,net1803);
INTERCONNECT SplitCLK_4_764_SplitCLK_6_762(net1804_c1,net1804);
INTERCONNECT SplitCLK_4_764_SplitCLK_6_763(net1805_c1,net1805);
INTERCONNECT SplitCLK_6_763_SplitCLK_2_1516(net1806_c1,net1806);
INTERCONNECT SplitCLK_6_763_SplitCLK_4_1535(net1807_c1,net1807);
INTERCONNECT SplitCLK_6_762_SplitCLK_2_1183(net1808_c1,net1808);
INTERCONNECT SplitCLK_6_762_SplitCLK_4_1186(net1809_c1,net1809);
INTERCONNECT SplitCLK_0_761_SplitCLK_4_759(net1810_c1,net1810);
INTERCONNECT SplitCLK_0_761_SplitCLK_4_760(net1811_c1,net1811);
INTERCONNECT SplitCLK_4_760_SplitCLK_2_1050(net1812_c1,net1812);
INTERCONNECT SplitCLK_4_760_SplitCLK_4_1067(net1813_c1,net1813);
INTERCONNECT SplitCLK_4_759_SplitCLK_2_1264(net1814_c1,net1814);
INTERCONNECT SplitCLK_4_759_SplitCLK_4_1274(net1815_c1,net1815);
INTERCONNECT SplitCLK_6_758_SplitCLK_0_754(net1816_c1,net1816);
INTERCONNECT SplitCLK_6_758_SplitCLK_4_757(net1817_c1,net1817);
INTERCONNECT SplitCLK_4_757_SplitCLK_6_755(net1818_c1,net1818);
INTERCONNECT SplitCLK_4_757_SplitCLK_6_756(net1819_c1,net1819);
INTERCONNECT SplitCLK_6_756_SplitCLK_2_1085(net1820_c1,net1820);
INTERCONNECT SplitCLK_6_756_SplitCLK_4_1086(net1821_c1,net1821);
INTERCONNECT SplitCLK_6_755_SplitCLK_4_1483(net1822_c1,net1822);
INTERCONNECT SplitCLK_6_755_SplitCLK_2_1506(net1823_c1,net1823);
INTERCONNECT SplitCLK_0_754_SplitCLK_4_752(net1824_c1,net1824);
INTERCONNECT SplitCLK_0_754_SplitCLK_4_753(net1825_c1,net1825);
INTERCONNECT SplitCLK_4_753_SplitCLK_2_1119(net1826_c1,net1826);
INTERCONNECT SplitCLK_4_753_SplitCLK_4_1128(net1827_c1,net1827);
INTERCONNECT SplitCLK_4_752_SplitCLK_2_1453(net1828_c1,net1828);
INTERCONNECT SplitCLK_4_752_SplitCLK_2_1456(net1829_c1,net1829);
INTERCONNECT SplitCLK_6_751_SplitCLK_0_735(net1830_c1,net1830);
INTERCONNECT SplitCLK_6_751_SplitCLK_2_750(net1831_c1,net1831);
INTERCONNECT SplitCLK_2_750_SplitCLK_6_742(net1832_c1,net1832);
INTERCONNECT SplitCLK_2_750_SplitCLK_4_749(net1833_c1,net1833);
INTERCONNECT SplitCLK_4_749_SplitCLK_0_745(net1834_c1,net1834);
INTERCONNECT SplitCLK_4_749_SplitCLK_2_748(net1835_c1,net1835);
INTERCONNECT SplitCLK_2_748_SplitCLK_6_746(net1836_c1,net1836);
INTERCONNECT SplitCLK_2_748_SplitCLK_4_747(net1837_c1,net1837);
INTERCONNECT SplitCLK_4_747_SplitCLK_4_1055(net1838_c1,net1838);
INTERCONNECT SplitCLK_4_747_SplitCLK_2_1141(net1839_c1,net1839);
INTERCONNECT SplitCLK_6_746_SplitCLK_2_1255(net1840_c1,net1840);
INTERCONNECT SplitCLK_6_746_SplitCLK_4_1503(net1841_c1,net1841);
INTERCONNECT SplitCLK_0_745_SplitCLK_4_743(net1842_c1,net1842);
INTERCONNECT SplitCLK_0_745_SplitCLK_4_744(net1843_c1,net1843);
INTERCONNECT SplitCLK_4_744_SplitCLK_2_1403(net1844_c1,net1844);
INTERCONNECT SplitCLK_4_744_SplitCLK_4_1465(net1845_c1,net1845);
INTERCONNECT SplitCLK_4_743_SplitCLK_4_1426(net1846_c1,net1846);
INTERCONNECT SplitCLK_4_743_SplitCLK_2_1479(net1847_c1,net1847);
INTERCONNECT SplitCLK_6_742_SplitCLK_4_738(net1848_c1,net1848);
INTERCONNECT SplitCLK_6_742_SplitCLK_6_741(net1849_c1,net1849);
INTERCONNECT SplitCLK_6_741_SplitCLK_6_739(net1850_c1,net1850);
INTERCONNECT SplitCLK_6_741_SplitCLK_4_740(net1851_c1,net1851);
INTERCONNECT SplitCLK_4_740_SplitCLK_2_1104(net1852_c1,net1852);
INTERCONNECT SplitCLK_4_740_SplitCLK_4_1355(net1853_c1,net1853);
INTERCONNECT SplitCLK_6_739_SplitCLK_4_1245(net1854_c1,net1854);
INTERCONNECT SplitCLK_6_739_SplitCLK_2_1541(net1855_c1,net1855);
INTERCONNECT SplitCLK_4_738_SplitCLK_6_736(net1856_c1,net1856);
INTERCONNECT SplitCLK_4_738_SplitCLK_0_737(net1857_c1,net1857);
INTERCONNECT SplitCLK_0_737_SplitCLK_4_1176(net1858_c1,net1858);
INTERCONNECT SplitCLK_0_737_SplitCLK_2_1262(net1859_c1,net1859);
INTERCONNECT SplitCLK_6_736_SplitCLK_4_1168(net1860_c1,net1860);
INTERCONNECT SplitCLK_6_736_SplitCLK_2_1344(net1861_c1,net1861);
INTERCONNECT SplitCLK_0_735_SplitCLK_6_727(net1862_c1,net1862);
INTERCONNECT SplitCLK_0_735_SplitCLK_4_734(net1863_c1,net1863);
INTERCONNECT SplitCLK_4_734_SplitCLK_4_730(net1864_c1,net1864);
INTERCONNECT SplitCLK_4_734_SplitCLK_2_733(net1865_c1,net1865);
INTERCONNECT SplitCLK_2_733_SplitCLK_2_731(net1866_c1,net1866);
INTERCONNECT SplitCLK_2_733_SplitCLK_4_732(net1867_c1,net1867);
INTERCONNECT SplitCLK_4_732_SplitCLK_4_1410(net1868_c1,net1868);
INTERCONNECT SplitCLK_4_732_SplitCLK_2_1449(net1869_c1,net1869);
INTERCONNECT SplitCLK_2_731_SplitCLK_2_1216(net1870_c1,net1870);
INTERCONNECT SplitCLK_2_731_SplitCLK_4_1409(net1871_c1,net1871);
INTERCONNECT SplitCLK_4_730_SplitCLK_0_728(net1872_c1,net1872);
INTERCONNECT SplitCLK_4_730_SplitCLK_4_729(net1873_c1,net1873);
INTERCONNECT SplitCLK_4_729_SplitCLK_2_1383(net1874_c1,net1874);
INTERCONNECT SplitCLK_4_729_SplitCLK_4_1432(net1875_c1,net1875);
INTERCONNECT SplitCLK_0_728_SplitCLK_4_1361(net1876_c1,net1876);
INTERCONNECT SplitCLK_0_728_SplitCLK_4_1401(net1877_c1,net1877);
INTERCONNECT SplitCLK_6_727_SplitCLK_4_723(net1878_c1,net1878);
INTERCONNECT SplitCLK_6_727_SplitCLK_6_726(net1879_c1,net1879);
INTERCONNECT SplitCLK_6_726_SplitCLK_6_724(net1880_c1,net1880);
INTERCONNECT SplitCLK_6_726_SplitCLK_4_725(net1881_c1,net1881);
INTERCONNECT SplitCLK_4_725_SplitCLK_4_1117(net1882_c1,net1882);
INTERCONNECT SplitCLK_4_725_SplitCLK_2_1241(net1883_c1,net1883);
INTERCONNECT SplitCLK_6_724_SplitCLK_2_1294(net1884_c1,net1884);
INTERCONNECT SplitCLK_6_724_SplitCLK_4_1308(net1885_c1,net1885);
INTERCONNECT SplitCLK_4_723_SplitCLK_4_721(net1886_c1,net1886);
INTERCONNECT SplitCLK_4_723_SplitCLK_4_722(net1887_c1,net1887);
INTERCONNECT SplitCLK_4_722_SplitCLK_4_1377(net1888_c1,net1888);
INTERCONNECT SplitCLK_4_722_SplitCLK_2_1384(net1889_c1,net1889);
INTERCONNECT SplitCLK_4_721_SplitCLK_2_1431(net1890_c1,net1890);
INTERCONNECT SplitCLK_4_721_SplitCLK_4_720(net1891_c1,net1891);
INTERCONNECT SplitCLK_4_720_OR2T_79_n80(net1892_c1,net1892);
INTERCONNECT SplitCLK_4_720_DFFT_236__FPB_n1416(net1893_c1,net1893);
INTERCONNECT SplitCLK_0_719_SplitCLK_6_686(net1894_c1,net1894);
INTERCONNECT SplitCLK_0_719_SplitCLK_4_718(net1895_c1,net1895);
INTERCONNECT SplitCLK_4_718_SplitCLK_0_702(net1896_c1,net1896);
INTERCONNECT SplitCLK_4_718_SplitCLK_4_717(net1897_c1,net1897);
INTERCONNECT SplitCLK_4_717_SplitCLK_6_709(net1898_c1,net1898);
INTERCONNECT SplitCLK_4_717_SplitCLK_4_716(net1899_c1,net1899);
INTERCONNECT SplitCLK_4_716_SplitCLK_0_712(net1900_c1,net1900);
INTERCONNECT SplitCLK_4_716_SplitCLK_4_715(net1901_c1,net1901);
INTERCONNECT SplitCLK_4_715_SplitCLK_6_713(net1902_c1,net1902);
INTERCONNECT SplitCLK_4_715_SplitCLK_6_714(net1903_c1,net1903);
INTERCONNECT SplitCLK_6_714_SplitCLK_2_1079(net1904_c1,net1904);
INTERCONNECT SplitCLK_6_714_SplitCLK_4_1444(net1905_c1,net1905);
INTERCONNECT SplitCLK_6_713_SplitCLK_2_1285(net1906_c1,net1906);
INTERCONNECT SplitCLK_6_713_SplitCLK_4_1301(net1907_c1,net1907);
INTERCONNECT SplitCLK_0_712_SplitCLK_4_710(net1908_c1,net1908);
INTERCONNECT SplitCLK_0_712_SplitCLK_4_711(net1909_c1,net1909);
INTERCONNECT SplitCLK_4_711_SplitCLK_2_1474(net1910_c1,net1910);
INTERCONNECT SplitCLK_4_711_SplitCLK_4_1497(net1911_c1,net1911);
INTERCONNECT SplitCLK_4_710_SplitCLK_2_1315(net1912_c1,net1912);
INTERCONNECT SplitCLK_4_710_SplitCLK_4_1353(net1913_c1,net1913);
INTERCONNECT SplitCLK_6_709_SplitCLK_0_705(net1914_c1,net1914);
INTERCONNECT SplitCLK_6_709_SplitCLK_2_708(net1915_c1,net1915);
INTERCONNECT SplitCLK_2_708_SplitCLK_6_706(net1916_c1,net1916);
INTERCONNECT SplitCLK_2_708_SplitCLK_4_707(net1917_c1,net1917);
INTERCONNECT SplitCLK_4_707_SplitCLK_2_1137(net1918_c1,net1918);
INTERCONNECT SplitCLK_4_707_SplitCLK_4_1396(net1919_c1,net1919);
INTERCONNECT SplitCLK_6_706_SplitCLK_2_1142(net1920_c1,net1920);
INTERCONNECT SplitCLK_6_706_SplitCLK_4_1146(net1921_c1,net1921);
INTERCONNECT SplitCLK_0_705_SplitCLK_4_703(net1922_c1,net1922);
INTERCONNECT SplitCLK_0_705_SplitCLK_4_704(net1923_c1,net1923);
INTERCONNECT SplitCLK_4_704_SplitCLK_4_1268(net1924_c1,net1924);
INTERCONNECT SplitCLK_4_704_SplitCLK_2_1375(net1925_c1,net1925);
INTERCONNECT SplitCLK_4_703_SplitCLK_2_1114(net1926_c1,net1926);
INTERCONNECT SplitCLK_4_703_SplitCLK_4_1305(net1927_c1,net1927);
INTERCONNECT SplitCLK_0_702_SplitCLK_4_694(net1928_c1,net1928);
INTERCONNECT SplitCLK_0_702_SplitCLK_4_701(net1929_c1,net1929);
INTERCONNECT SplitCLK_4_701_SplitCLK_4_697(net1930_c1,net1930);
INTERCONNECT SplitCLK_4_701_SplitCLK_2_700(net1931_c1,net1931);
INTERCONNECT SplitCLK_2_700_SplitCLK_6_698(net1932_c1,net1932);
INTERCONNECT SplitCLK_2_700_SplitCLK_4_699(net1933_c1,net1933);
INTERCONNECT SplitCLK_4_699_SplitCLK_2_1515(net1934_c1,net1934);
INTERCONNECT SplitCLK_4_699_SplitCLK_4_1534(net1935_c1,net1935);
INTERCONNECT SplitCLK_6_698_SplitCLK_2_1278(net1936_c1,net1936);
INTERCONNECT SplitCLK_6_698_SplitCLK_4_1334(net1937_c1,net1937);
INTERCONNECT SplitCLK_4_697_SplitCLK_0_695(net1938_c1,net1938);
INTERCONNECT SplitCLK_4_697_SplitCLK_4_696(net1939_c1,net1939);
INTERCONNECT SplitCLK_4_696_SplitCLK_4_1049(net1940_c1,net1940);
INTERCONNECT SplitCLK_4_696_SplitCLK_2_1066(net1941_c1,net1941);
INTERCONNECT SplitCLK_0_695_SplitCLK_4_1078(net1942_c1,net1942);
INTERCONNECT SplitCLK_0_695_SplitCLK_4_1090(net1943_c1,net1943);
INTERCONNECT SplitCLK_4_694_SplitCLK_4_690(net1944_c1,net1944);
INTERCONNECT SplitCLK_4_694_SplitCLK_6_693(net1945_c1,net1945);
INTERCONNECT SplitCLK_6_693_SplitCLK_6_691(net1946_c1,net1946);
INTERCONNECT SplitCLK_6_693_SplitCLK_2_692(net1947_c1,net1947);
INTERCONNECT SplitCLK_2_692_SplitCLK_4_1291(net1948_c1,net1948);
INTERCONNECT SplitCLK_2_692_SplitCLK_2_1321(net1949_c1,net1949);
INTERCONNECT SplitCLK_6_691_SplitCLK_4_1402(net1950_c1,net1950);
INTERCONNECT SplitCLK_6_691_SplitCLK_2_1425(net1951_c1,net1951);
INTERCONNECT SplitCLK_4_690_SplitCLK_0_688(net1952_c1,net1952);
INTERCONNECT SplitCLK_4_690_SplitCLK_2_689(net1953_c1,net1953);
INTERCONNECT SplitCLK_2_689_SplitCLK_2_1103(net1954_c1,net1954);
INTERCONNECT SplitCLK_2_689_SplitCLK_4_1123(net1955_c1,net1955);
INTERCONNECT SplitCLK_0_688_SplitCLK_2_1130(net1956_c1,net1956);
INTERCONNECT SplitCLK_0_688_SplitCLK_4_687(net1957_c1,net1957);
INTERCONNECT SplitCLK_4_687_XOR2T_134_R0(net1958_c1,net1958);
INTERCONNECT SplitCLK_4_687_AND2T_135_n136(net1959_c1,net1959);
INTERCONNECT SplitCLK_6_686_SplitCLK_0_670(net1960_c1,net1960);
INTERCONNECT SplitCLK_6_686_SplitCLK_2_685(net1961_c1,net1961);
INTERCONNECT SplitCLK_2_685_SplitCLK_6_677(net1962_c1,net1962);
INTERCONNECT SplitCLK_2_685_SplitCLK_4_684(net1963_c1,net1963);
INTERCONNECT SplitCLK_4_684_SplitCLK_4_680(net1964_c1,net1964);
INTERCONNECT SplitCLK_4_684_SplitCLK_2_683(net1965_c1,net1965);
INTERCONNECT SplitCLK_2_683_SplitCLK_0_681(net1966_c1,net1966);
INTERCONNECT SplitCLK_2_683_SplitCLK_2_682(net1967_c1,net1967);
INTERCONNECT SplitCLK_2_682_SplitCLK_4_1486(net1968_c1,net1968);
INTERCONNECT SplitCLK_2_682_SplitCLK_2_1527(net1969_c1,net1969);
INTERCONNECT SplitCLK_0_681_SplitCLK_2_1424(net1970_c1,net1970);
INTERCONNECT SplitCLK_0_681_SplitCLK_4_1509(net1971_c1,net1971);
INTERCONNECT SplitCLK_4_680_SplitCLK_6_678(net1972_c1,net1972);
INTERCONNECT SplitCLK_4_680_SplitCLK_4_679(net1973_c1,net1973);
INTERCONNECT SplitCLK_4_679_SplitCLK_2_1336(net1974_c1,net1974);
INTERCONNECT SplitCLK_4_679_SplitCLK_4_1356(net1975_c1,net1975);
INTERCONNECT SplitCLK_6_678_SplitCLK_4_1500(net1976_c1,net1976);
INTERCONNECT SplitCLK_6_678_SplitCLK_2_1518(net1977_c1,net1977);
INTERCONNECT SplitCLK_6_677_SplitCLK_4_673(net1978_c1,net1978);
INTERCONNECT SplitCLK_6_677_SplitCLK_6_676(net1979_c1,net1979);
INTERCONNECT SplitCLK_6_676_SplitCLK_6_674(net1980_c1,net1980);
INTERCONNECT SplitCLK_6_676_SplitCLK_4_675(net1981_c1,net1981);
INTERCONNECT SplitCLK_4_675_SplitCLK_4_1107(net1982_c1,net1982);
INTERCONNECT SplitCLK_4_675_SplitCLK_2_1446(net1983_c1,net1983);
INTERCONNECT SplitCLK_6_674_SplitCLK_4_1214(net1984_c1,net1984);
INTERCONNECT SplitCLK_6_674_SplitCLK_2_1343(net1985_c1,net1985);
INTERCONNECT SplitCLK_4_673_SplitCLK_0_671(net1986_c1,net1986);
INTERCONNECT SplitCLK_4_673_SplitCLK_4_672(net1987_c1,net1987);
INTERCONNECT SplitCLK_4_672_SplitCLK_4_1110(net1988_c1,net1988);
INTERCONNECT SplitCLK_4_672_SplitCLK_2_1476(net1989_c1,net1989);
INTERCONNECT SplitCLK_0_671_SplitCLK_2_1177(net1990_c1,net1990);
INTERCONNECT SplitCLK_0_671_SplitCLK_4_1499(net1991_c1,net1991);
INTERCONNECT SplitCLK_0_670_SplitCLK_6_662(net1992_c1,net1992);
INTERCONNECT SplitCLK_0_670_SplitCLK_4_669(net1993_c1,net1993);
INTERCONNECT SplitCLK_4_669_SplitCLK_4_665(net1994_c1,net1994);
INTERCONNECT SplitCLK_4_669_SplitCLK_6_668(net1995_c1,net1995);
INTERCONNECT SplitCLK_6_668_SplitCLK_0_666(net1996_c1,net1996);
INTERCONNECT SplitCLK_6_668_SplitCLK_0_667(net1997_c1,net1997);
INTERCONNECT SplitCLK_0_667_SplitCLK_4_1378(net1998_c1,net1998);
INTERCONNECT SplitCLK_0_667_SplitCLK_2_1477(net1999_c1,net1999);
INTERCONNECT SplitCLK_0_666_SplitCLK_2_1190(net2000_c1,net2000);
INTERCONNECT SplitCLK_0_666_SplitCLK_4_1447(net2001_c1,net2001);
INTERCONNECT SplitCLK_4_665_SplitCLK_0_663(net2002_c1,net2002);
INTERCONNECT SplitCLK_4_665_SplitCLK_4_664(net2003_c1,net2003);
INTERCONNECT SplitCLK_4_664_SplitCLK_4_1088(net2004_c1,net2004);
INTERCONNECT SplitCLK_4_664_SplitCLK_2_1121(net2005_c1,net2005);
INTERCONNECT SplitCLK_0_663_SplitCLK_4_1076(net2006_c1,net2006);
INTERCONNECT SplitCLK_0_663_SplitCLK_2_1536(net2007_c1,net2007);
INTERCONNECT SplitCLK_6_662_SplitCLK_0_658(net2008_c1,net2008);
INTERCONNECT SplitCLK_6_662_SplitCLK_2_661(net2009_c1,net2009);
INTERCONNECT SplitCLK_2_661_SplitCLK_0_659(net2010_c1,net2010);
INTERCONNECT SplitCLK_2_661_SplitCLK_6_660(net2011_c1,net2011);
INTERCONNECT SplitCLK_6_660_SplitCLK_4_1064(net2012_c1,net2012);
INTERCONNECT SplitCLK_6_660_SplitCLK_2_1517(net2013_c1,net2013);
INTERCONNECT SplitCLK_0_659_SplitCLK_4_1048(net2014_c1,net2014);
INTERCONNECT SplitCLK_0_659_SplitCLK_2_1242(net2015_c1,net2015);
INTERCONNECT SplitCLK_0_658_SplitCLK_6_656(net2016_c1,net2016);
INTERCONNECT SplitCLK_0_658_SplitCLK_4_657(net2017_c1,net2017);
INTERCONNECT SplitCLK_4_657_SplitCLK_2_1051(net2018_c1,net2018);
INTERCONNECT SplitCLK_4_657_SplitCLK_4_1400(net2019_c1,net2019);
INTERCONNECT SplitCLK_6_656_SplitCLK_2_1306(net2020_c1,net2020);
INTERCONNECT SplitCLK_6_656_SplitCLK_4_655(net2021_c1,net2021);
INTERCONNECT SplitCLK_4_655_DFFT_469__FPB_n1649(net2022_c1,net2022);
INTERCONNECT SplitCLK_4_655_DFFT_470__FPB_n1650(net2023_c1,net2023);
INTERCONNECT SplitCLK_6_654_SplitCLK_0_589(net2024_c1,net2024);
INTERCONNECT SplitCLK_6_654_SplitCLK_2_653(net2025_c1,net2025);
INTERCONNECT SplitCLK_2_653_SplitCLK_6_621(net2026_c1,net2026);
INTERCONNECT SplitCLK_2_653_SplitCLK_4_652(net2027_c1,net2027);
INTERCONNECT SplitCLK_4_652_SplitCLK_0_636(net2028_c1,net2028);
INTERCONNECT SplitCLK_4_652_SplitCLK_2_651(net2029_c1,net2029);
INTERCONNECT SplitCLK_2_651_SplitCLK_6_643(net2030_c1,net2030);
INTERCONNECT SplitCLK_2_651_SplitCLK_4_650(net2031_c1,net2031);
INTERCONNECT SplitCLK_4_650_SplitCLK_0_646(net2032_c1,net2032);
INTERCONNECT SplitCLK_4_650_SplitCLK_4_649(net2033_c1,net2033);
INTERCONNECT SplitCLK_4_649_SplitCLK_6_647(net2034_c1,net2034);
INTERCONNECT SplitCLK_4_649_SplitCLK_6_648(net2035_c1,net2035);
INTERCONNECT SplitCLK_6_648_SplitCLK_2_1450(net2036_c1,net2036);
INTERCONNECT SplitCLK_6_648_SplitCLK_4_1480(net2037_c1,net2037);
INTERCONNECT SplitCLK_6_647_SplitCLK_2_1357(net2038_c1,net2038);
INTERCONNECT SplitCLK_6_647_SplitCLK_4_1523(net2039_c1,net2039);
INTERCONNECT SplitCLK_0_646_SplitCLK_4_644(net2040_c1,net2040);
INTERCONNECT SplitCLK_0_646_SplitCLK_4_645(net2041_c1,net2041);
INTERCONNECT SplitCLK_4_645_SplitCLK_4_1427(net2042_c1,net2042);
INTERCONNECT SplitCLK_4_645_SplitCLK_2_1504(net2043_c1,net2043);
INTERCONNECT SplitCLK_4_644_SplitCLK_4_1106(net2044_c1,net2044);
INTERCONNECT SplitCLK_4_644_SplitCLK_2_1467(net2045_c1,net2045);
INTERCONNECT SplitCLK_6_643_SplitCLK_4_639(net2046_c1,net2046);
INTERCONNECT SplitCLK_6_643_SplitCLK_6_642(net2047_c1,net2047);
INTERCONNECT SplitCLK_6_642_SplitCLK_4_640(net2048_c1,net2048);
INTERCONNECT SplitCLK_6_642_SplitCLK_4_641(net2049_c1,net2049);
INTERCONNECT SplitCLK_4_641_SplitCLK_4_1163(net2050_c1,net2050);
INTERCONNECT SplitCLK_4_641_SplitCLK_2_1436(net2051_c1,net2051);
INTERCONNECT SplitCLK_4_640_SplitCLK_2_1235(net2052_c1,net2052);
INTERCONNECT SplitCLK_4_640_SplitCLK_2_1250(net2053_c1,net2053);
INTERCONNECT SplitCLK_4_639_SplitCLK_6_637(net2054_c1,net2054);
INTERCONNECT SplitCLK_4_639_SplitCLK_2_638(net2055_c1,net2055);
INTERCONNECT SplitCLK_2_638_SplitCLK_4_1174(net2056_c1,net2056);
INTERCONNECT SplitCLK_2_638_SplitCLK_2_1237(net2057_c1,net2057);
INTERCONNECT SplitCLK_6_637_SplitCLK_4_1184(net2058_c1,net2058);
INTERCONNECT SplitCLK_6_637_SplitCLK_2_1542(net2059_c1,net2059);
INTERCONNECT SplitCLK_0_636_SplitCLK_6_628(net2060_c1,net2060);
INTERCONNECT SplitCLK_0_636_SplitCLK_4_635(net2061_c1,net2061);
INTERCONNECT SplitCLK_4_635_SplitCLK_4_631(net2062_c1,net2062);
INTERCONNECT SplitCLK_4_635_SplitCLK_2_634(net2063_c1,net2063);
INTERCONNECT SplitCLK_2_634_SplitCLK_0_632(net2064_c1,net2064);
INTERCONNECT SplitCLK_2_634_SplitCLK_4_633(net2065_c1,net2065);
INTERCONNECT SplitCLK_4_633_SplitCLK_2_1380(net2066_c1,net2066);
INTERCONNECT SplitCLK_4_633_SplitCLK_2_1405(net2067_c1,net2067);
INTERCONNECT SplitCLK_0_632_SplitCLK_2_1293(net2068_c1,net2068);
INTERCONNECT SplitCLK_0_632_SplitCLK_4_1358(net2069_c1,net2069);
INTERCONNECT SplitCLK_4_631_SplitCLK_0_629(net2070_c1,net2070);
INTERCONNECT SplitCLK_4_631_SplitCLK_4_630(net2071_c1,net2071);
INTERCONNECT SplitCLK_4_630_SplitCLK_4_1213(net2072_c1,net2072);
INTERCONNECT SplitCLK_4_630_SplitCLK_2_1362(net2073_c1,net2073);
INTERCONNECT SplitCLK_0_629_SplitCLK_2_1337(net2074_c1,net2074);
INTERCONNECT SplitCLK_0_629_SplitCLK_4_1340(net2075_c1,net2075);
INTERCONNECT SplitCLK_6_628_SplitCLK_4_624(net2076_c1,net2076);
INTERCONNECT SplitCLK_6_628_SplitCLK_6_627(net2077_c1,net2077);
INTERCONNECT SplitCLK_6_627_SplitCLK_6_625(net2078_c1,net2078);
INTERCONNECT SplitCLK_6_627_SplitCLK_4_626(net2079_c1,net2079);
INTERCONNECT SplitCLK_4_626_SplitCLK_2_1172(net2080_c1,net2080);
INTERCONNECT SplitCLK_4_626_SplitCLK_4_1279(net2081_c1,net2081);
INTERCONNECT SplitCLK_6_625_SplitCLK_4_1217(net2082_c1,net2082);
INTERCONNECT SplitCLK_6_625_SplitCLK_2_1234(net2083_c1,net2083);
INTERCONNECT SplitCLK_4_624_SplitCLK_0_622(net2084_c1,net2084);
INTERCONNECT SplitCLK_4_624_SplitCLK_4_623(net2085_c1,net2085);
INTERCONNECT SplitCLK_4_623_SplitCLK_2_1269(net2086_c1,net2086);
INTERCONNECT SplitCLK_4_623_SplitCLK_4_1387(net2087_c1,net2087);
INTERCONNECT SplitCLK_0_622_SplitCLK_4_1171(net2088_c1,net2088);
INTERCONNECT SplitCLK_0_622_SplitCLK_2_1227(net2089_c1,net2089);
INTERCONNECT SplitCLK_6_621_SplitCLK_0_605(net2090_c1,net2090);
INTERCONNECT SplitCLK_6_621_SplitCLK_6_620(net2091_c1,net2091);
INTERCONNECT SplitCLK_6_620_SplitCLK_6_612(net2092_c1,net2092);
INTERCONNECT SplitCLK_6_620_SplitCLK_4_619(net2093_c1,net2093);
INTERCONNECT SplitCLK_4_619_SplitCLK_4_615(net2094_c1,net2094);
INTERCONNECT SplitCLK_4_619_SplitCLK_6_618(net2095_c1,net2095);
INTERCONNECT SplitCLK_6_618_SplitCLK_6_616(net2096_c1,net2096);
INTERCONNECT SplitCLK_6_618_SplitCLK_4_617(net2097_c1,net2097);
INTERCONNECT SplitCLK_4_617_SplitCLK_2_1154(net2098_c1,net2098);
INTERCONNECT SplitCLK_4_617_SplitCLK_4_1202(net2099_c1,net2099);
INTERCONNECT SplitCLK_6_616_SplitCLK_4_1209(net2100_c1,net2100);
INTERCONNECT SplitCLK_6_616_SplitCLK_2_1488(net2101_c1,net2101);
INTERCONNECT SplitCLK_4_615_SplitCLK_2_613(net2102_c1,net2102);
INTERCONNECT SplitCLK_4_615_SplitCLK_4_614(net2103_c1,net2103);
INTERCONNECT SplitCLK_4_614_SplitCLK_4_1169(net2104_c1,net2104);
INTERCONNECT SplitCLK_4_614_SplitCLK_4_1459(net2105_c1,net2105);
INTERCONNECT SplitCLK_2_613_SplitCLK_2_1205(net2106_c1,net2106);
INTERCONNECT SplitCLK_2_613_SplitCLK_2_1211(net2107_c1,net2107);
INTERCONNECT SplitCLK_6_612_SplitCLK_0_608(net2108_c1,net2108);
INTERCONNECT SplitCLK_6_612_SplitCLK_6_611(net2109_c1,net2109);
INTERCONNECT SplitCLK_6_611_SplitCLK_6_609(net2110_c1,net2110);
INTERCONNECT SplitCLK_6_611_SplitCLK_4_610(net2111_c1,net2111);
INTERCONNECT SplitCLK_4_610_SplitCLK_4_1283(net2112_c1,net2112);
INTERCONNECT SplitCLK_4_610_SplitCLK_2_1421(net2113_c1,net2113);
INTERCONNECT SplitCLK_6_609_SplitCLK_2_1473(net2114_c1,net2114);
INTERCONNECT SplitCLK_6_609_SplitCLK_4_1495(net2115_c1,net2115);
INTERCONNECT SplitCLK_0_608_SplitCLK_6_606(net2116_c1,net2116);
INTERCONNECT SplitCLK_0_608_SplitCLK_0_607(net2117_c1,net2117);
INTERCONNECT SplitCLK_0_607_SplitCLK_2_1298(net2118_c1,net2118);
INTERCONNECT SplitCLK_0_607_SplitCLK_4_1420(net2119_c1,net2119);
INTERCONNECT SplitCLK_6_606_SplitCLK_2_1514(net2120_c1,net2120);
INTERCONNECT SplitCLK_6_606_SplitCLK_4_1532(net2121_c1,net2121);
INTERCONNECT SplitCLK_0_605_SplitCLK_6_597(net2122_c1,net2122);
INTERCONNECT SplitCLK_0_605_SplitCLK_4_604(net2123_c1,net2123);
INTERCONNECT SplitCLK_4_604_SplitCLK_0_600(net2124_c1,net2124);
INTERCONNECT SplitCLK_4_604_SplitCLK_4_603(net2125_c1,net2125);
INTERCONNECT SplitCLK_4_603_SplitCLK_6_601(net2126_c1,net2126);
INTERCONNECT SplitCLK_4_603_SplitCLK_6_602(net2127_c1,net2127);
INTERCONNECT SplitCLK_6_602_SplitCLK_4_1098(net2128_c1,net2128);
INTERCONNECT SplitCLK_6_602_SplitCLK_2_1164(net2129_c1,net2129);
INTERCONNECT SplitCLK_6_601_SplitCLK_2_1165(net2130_c1,net2130);
INTERCONNECT SplitCLK_6_601_SplitCLK_2_1460(net2131_c1,net2131);
INTERCONNECT SplitCLK_0_600_SplitCLK_4_598(net2132_c1,net2132);
INTERCONNECT SplitCLK_0_600_SplitCLK_4_599(net2133_c1,net2133);
INTERCONNECT SplitCLK_4_599_SplitCLK_4_1153(net2134_c1,net2134);
INTERCONNECT SplitCLK_4_599_SplitCLK_2_1222(net2135_c1,net2135);
INTERCONNECT SplitCLK_4_598_SplitCLK_2_1188(net2136_c1,net2136);
INTERCONNECT SplitCLK_4_598_SplitCLK_4_1347(net2137_c1,net2137);
INTERCONNECT SplitCLK_6_597_SplitCLK_0_593(net2138_c1,net2138);
INTERCONNECT SplitCLK_6_597_SplitCLK_6_596(net2139_c1,net2139);
INTERCONNECT SplitCLK_6_596_SplitCLK_6_594(net2140_c1,net2140);
INTERCONNECT SplitCLK_6_596_SplitCLK_4_595(net2141_c1,net2141);
INTERCONNECT SplitCLK_4_595_SplitCLK_2_1443(net2142_c1,net2142);
INTERCONNECT SplitCLK_4_595_SplitCLK_4_1470(net2143_c1,net2143);
INTERCONNECT SplitCLK_6_594_SplitCLK_4_1074(net2144_c1,net2144);
INTERCONNECT SplitCLK_6_594_SplitCLK_2_1136(net2145_c1,net2145);
INTERCONNECT SplitCLK_0_593_SplitCLK_6_591(net2146_c1,net2146);
INTERCONNECT SplitCLK_0_593_SplitCLK_4_592(net2147_c1,net2147);
INTERCONNECT SplitCLK_4_592_SplitCLK_4_1166(net2148_c1,net2148);
INTERCONNECT SplitCLK_4_592_SplitCLK_2_1212(net2149_c1,net2149);
INTERCONNECT SplitCLK_6_591_SplitCLK_2_1062(net2150_c1,net2150);
INTERCONNECT SplitCLK_6_591_SplitCLK_4_590(net2151_c1,net2151);
INTERCONNECT SplitCLK_4_590_XOR2T_47_n48(net2152_c1,net2152);
INTERCONNECT SplitCLK_4_590_DFFT_143__FPB_n144(net2153_c1,net2153);
INTERCONNECT SplitCLK_0_589_SplitCLK_6_556(net2154_c1,net2154);
INTERCONNECT SplitCLK_0_589_SplitCLK_4_588(net2155_c1,net2155);
INTERCONNECT SplitCLK_4_588_SplitCLK_4_572(net2156_c1,net2156);
INTERCONNECT SplitCLK_4_588_SplitCLK_2_587(net2157_c1,net2157);
INTERCONNECT SplitCLK_2_587_SplitCLK_2_579(net2158_c1,net2158);
INTERCONNECT SplitCLK_2_587_SplitCLK_4_586(net2159_c1,net2159);
INTERCONNECT SplitCLK_4_586_SplitCLK_0_582(net2160_c1,net2160);
INTERCONNECT SplitCLK_4_586_SplitCLK_2_585(net2161_c1,net2161);
INTERCONNECT SplitCLK_2_585_SplitCLK_6_583(net2162_c1,net2162);
INTERCONNECT SplitCLK_2_585_SplitCLK_4_584(net2163_c1,net2163);
INTERCONNECT SplitCLK_4_584_SplitCLK_2_1322(net2164_c1,net2164);
INTERCONNECT SplitCLK_4_584_SplitCLK_4_1487(net2165_c1,net2165);
INTERCONNECT SplitCLK_6_583_SplitCLK_2_1319(net2166_c1,net2166);
INTERCONNECT SplitCLK_6_583_SplitCLK_4_1363(net2167_c1,net2167);
INTERCONNECT SplitCLK_0_582_SplitCLK_6_580(net2168_c1,net2168);
INTERCONNECT SplitCLK_0_582_SplitCLK_4_581(net2169_c1,net2169);
INTERCONNECT SplitCLK_4_581_SplitCLK_4_1412(net2170_c1,net2170);
INTERCONNECT SplitCLK_4_581_SplitCLK_2_1457(net2171_c1,net2171);
INTERCONNECT SplitCLK_6_580_SplitCLK_2_1385(net2172_c1,net2172);
INTERCONNECT SplitCLK_6_580_SplitCLK_4_1411(net2173_c1,net2173);
INTERCONNECT SplitCLK_2_579_SplitCLK_4_575(net2174_c1,net2174);
INTERCONNECT SplitCLK_2_579_SplitCLK_2_578(net2175_c1,net2175);
INTERCONNECT SplitCLK_2_578_SplitCLK_6_576(net2176_c1,net2176);
INTERCONNECT SplitCLK_2_578_SplitCLK_4_577(net2177_c1,net2177);
INTERCONNECT SplitCLK_4_577_SplitCLK_4_1452(net2178_c1,net2178);
INTERCONNECT SplitCLK_4_577_SplitCLK_2_1482(net2179_c1,net2179);
INTERCONNECT SplitCLK_6_576_SplitCLK_2_1231(net2180_c1,net2180);
INTERCONNECT SplitCLK_6_576_SplitCLK_4_1239(net2181_c1,net2181);
INTERCONNECT SplitCLK_4_575_SplitCLK_6_573(net2182_c1,net2182);
INTERCONNECT SplitCLK_4_575_SplitCLK_4_574(net2183_c1,net2183);
INTERCONNECT SplitCLK_4_574_SplitCLK_2_1428(net2184_c1,net2184);
INTERCONNECT SplitCLK_4_574_SplitCLK_4_1433(net2185_c1,net2185);
INTERCONNECT SplitCLK_6_573_SplitCLK_2_1381(net2186_c1,net2186);
INTERCONNECT SplitCLK_6_573_SplitCLK_4_1406(net2187_c1,net2187);
INTERCONNECT SplitCLK_4_572_SplitCLK_6_564(net2188_c1,net2188);
INTERCONNECT SplitCLK_4_572_SplitCLK_0_571(net2189_c1,net2189);
INTERCONNECT SplitCLK_0_571_SplitCLK_0_567(net2190_c1,net2190);
INTERCONNECT SplitCLK_0_571_SplitCLK_2_570(net2191_c1,net2191);
INTERCONNECT SplitCLK_2_570_SplitCLK_4_568(net2192_c1,net2192);
INTERCONNECT SplitCLK_2_570_SplitCLK_4_569(net2193_c1,net2193);
INTERCONNECT SplitCLK_4_569_SplitCLK_4_1292(net2194_c1,net2194);
INTERCONNECT SplitCLK_4_569_SplitCLK_2_1434(net2195_c1,net2195);
INTERCONNECT SplitCLK_4_568_SplitCLK_2_1089(net2196_c1,net2196);
INTERCONNECT SplitCLK_4_568_SplitCLK_2_1364(net2197_c1,net2197);
INTERCONNECT SplitCLK_0_567_SplitCLK_4_565(net2198_c1,net2198);
INTERCONNECT SplitCLK_0_567_SplitCLK_4_566(net2199_c1,net2199);
INTERCONNECT SplitCLK_4_566_SplitCLK_2_1122(net2200_c1,net2200);
INTERCONNECT SplitCLK_4_566_SplitCLK_4_1131(net2201_c1,net2201);
INTERCONNECT SplitCLK_4_565_SplitCLK_2_1065(net2202_c1,net2202);
INTERCONNECT SplitCLK_4_565_SplitCLK_4_1077(net2203_c1,net2203);
INTERCONNECT SplitCLK_6_564_SplitCLK_4_560(net2204_c1,net2204);
INTERCONNECT SplitCLK_6_564_SplitCLK_6_563(net2205_c1,net2205);
INTERCONNECT SplitCLK_6_563_SplitCLK_6_561(net2206_c1,net2206);
INTERCONNECT SplitCLK_6_563_SplitCLK_2_562(net2207_c1,net2207);
INTERCONNECT SplitCLK_2_562_SplitCLK_2_1324(net2208_c1,net2208);
INTERCONNECT SplitCLK_2_562_SplitCLK_4_1386(net2209_c1,net2209);
INTERCONNECT SplitCLK_6_561_SplitCLK_4_1307(net2210_c1,net2210);
INTERCONNECT SplitCLK_6_561_SplitCLK_2_1365(net2211_c1,net2211);
INTERCONNECT SplitCLK_4_560_SplitCLK_0_558(net2212_c1,net2212);
INTERCONNECT SplitCLK_4_560_SplitCLK_6_559(net2213_c1,net2213);
INTERCONNECT SplitCLK_6_559_SplitCLK_2_1342(net2214_c1,net2214);
INTERCONNECT SplitCLK_6_559_SplitCLK_4_1533(net2215_c1,net2215);
INTERCONNECT SplitCLK_0_558_SplitCLK_2_1496(net2216_c1,net2216);
INTERCONNECT SplitCLK_0_558_SplitCLK_4_557(net2217_c1,net2217);
INTERCONNECT SplitCLK_4_557_DFFT_463__FPB_n1643(net2218_c1,net2218);
INTERCONNECT SplitCLK_4_557_DFFT_461__FPB_n1641(net2219_c1,net2219);
INTERCONNECT SplitCLK_6_556_SplitCLK_0_540(net2220_c1,net2220);
INTERCONNECT SplitCLK_6_556_SplitCLK_2_555(net2221_c1,net2221);
INTERCONNECT SplitCLK_2_555_SplitCLK_6_547(net2222_c1,net2222);
INTERCONNECT SplitCLK_2_555_SplitCLK_4_554(net2223_c1,net2223);
INTERCONNECT SplitCLK_4_554_SplitCLK_4_550(net2224_c1,net2224);
INTERCONNECT SplitCLK_4_554_SplitCLK_6_553(net2225_c1,net2225);
INTERCONNECT SplitCLK_6_553_SplitCLK_6_551(net2226_c1,net2226);
INTERCONNECT SplitCLK_6_553_SplitCLK_4_552(net2227_c1,net2227);
INTERCONNECT SplitCLK_4_552_SplitCLK_2_1199(net2228_c1,net2228);
INTERCONNECT SplitCLK_4_552_SplitCLK_4_1369(net2229_c1,net2229);
INTERCONNECT SplitCLK_6_551_SplitCLK_4_1311(net2230_c1,net2230);
INTERCONNECT SplitCLK_6_551_SplitCLK_2_1328(net2231_c1,net2231);
INTERCONNECT SplitCLK_4_550_SplitCLK_6_548(net2232_c1,net2232);
INTERCONNECT SplitCLK_4_550_SplitCLK_4_549(net2233_c1,net2233);
INTERCONNECT SplitCLK_4_549_SplitCLK_2_1167(net2234_c1,net2234);
INTERCONNECT SplitCLK_4_549_SplitCLK_4_1471(net2235_c1,net2235);
INTERCONNECT SplitCLK_6_548_SplitCLK_2_1297(net2236_c1,net2236);
INTERCONNECT SplitCLK_6_548_SplitCLK_4_1510(net2237_c1,net2237);
INTERCONNECT SplitCLK_6_547_SplitCLK_4_543(net2238_c1,net2238);
INTERCONNECT SplitCLK_6_547_SplitCLK_6_546(net2239_c1,net2239);
INTERCONNECT SplitCLK_6_546_SplitCLK_6_544(net2240_c1,net2240);
INTERCONNECT SplitCLK_6_546_SplitCLK_6_545(net2241_c1,net2241);
INTERCONNECT SplitCLK_6_545_SplitCLK_4_1159(net2242_c1,net2242);
INTERCONNECT SplitCLK_6_545_SplitCLK_2_1312(net2243_c1,net2243);
INTERCONNECT SplitCLK_6_544_SplitCLK_2_1118(net2244_c1,net2244);
INTERCONNECT SplitCLK_6_544_SplitCLK_4_1240(net2245_c1,net2245);
INTERCONNECT SplitCLK_4_543_SplitCLK_6_541(net2246_c1,net2246);
INTERCONNECT SplitCLK_4_543_SplitCLK_4_542(net2247_c1,net2247);
INTERCONNECT SplitCLK_4_542_SplitCLK_4_1207(net2248_c1,net2248);
INTERCONNECT SplitCLK_4_542_SplitCLK_2_1329(net2249_c1,net2249);
INTERCONNECT SplitCLK_6_541_SplitCLK_2_1096(net2250_c1,net2250);
INTERCONNECT SplitCLK_6_541_SplitCLK_2_1203(net2251_c1,net2251);
INTERCONNECT SplitCLK_0_540_SplitCLK_6_532(net2252_c1,net2252);
INTERCONNECT SplitCLK_0_540_SplitCLK_4_539(net2253_c1,net2253);
INTERCONNECT SplitCLK_4_539_SplitCLK_4_535(net2254_c1,net2254);
INTERCONNECT SplitCLK_4_539_SplitCLK_6_538(net2255_c1,net2255);
INTERCONNECT SplitCLK_6_538_SplitCLK_4_536(net2256_c1,net2256);
INTERCONNECT SplitCLK_6_538_SplitCLK_2_537(net2257_c1,net2257);
INTERCONNECT SplitCLK_2_537_SplitCLK_4_1376(net2258_c1,net2258);
INTERCONNECT SplitCLK_2_537_SplitCLK_2_1528(net2259_c1,net2259);
INTERCONNECT SplitCLK_4_536_SplitCLK_2_1490(net2260_c1,net2260);
INTERCONNECT SplitCLK_4_536_SplitCLK_2_1545(net2261_c1,net2261);
INTERCONNECT SplitCLK_4_535_SplitCLK_0_533(net2262_c1,net2262);
INTERCONNECT SplitCLK_4_535_SplitCLK_6_534(net2263_c1,net2263);
INTERCONNECT SplitCLK_6_534_SplitCLK_4_1059(net2264_c1,net2264);
INTERCONNECT SplitCLK_6_534_SplitCLK_4_1099(net2265_c1,net2265);
INTERCONNECT SplitCLK_0_533_SplitCLK_4_1181(net2266_c1,net2266);
INTERCONNECT SplitCLK_0_533_SplitCLK_2_1232(net2267_c1,net2267);
INTERCONNECT SplitCLK_6_532_SplitCLK_4_528(net2268_c1,net2268);
INTERCONNECT SplitCLK_6_532_SplitCLK_2_531(net2269_c1,net2269);
INTERCONNECT SplitCLK_2_531_SplitCLK_6_529(net2270_c1,net2270);
INTERCONNECT SplitCLK_2_531_SplitCLK_4_530(net2271_c1,net2271);
INTERCONNECT SplitCLK_4_530_SplitCLK_2_1201(net2272_c1,net2272);
INTERCONNECT SplitCLK_4_530_SplitCLK_4_1326(net2273_c1,net2273);
INTERCONNECT SplitCLK_6_529_SplitCLK_2_1348(net2274_c1,net2274);
INTERCONNECT SplitCLK_6_529_SplitCLK_4_1388(net2275_c1,net2275);
INTERCONNECT SplitCLK_4_528_SplitCLK_6_526(net2276_c1,net2276);
INTERCONNECT SplitCLK_4_528_SplitCLK_2_527(net2277_c1,net2277);
INTERCONNECT SplitCLK_2_527_SplitCLK_2_1170(net2278_c1,net2278);
INTERCONNECT SplitCLK_2_527_SplitCLK_4_1366(net2279_c1,net2279);
INTERCONNECT SplitCLK_6_526_SplitCLK_2_1489(net2280_c1,net2280);
INTERCONNECT SplitCLK_6_526_SplitCLK_4_525(net2281_c1,net2281);
INTERCONNECT SplitCLK_4_525_DFFT_188__FPB_n1368(net2282_c1,net2282);
INTERCONNECT SplitCLK_4_525_DFFT_189__FPB_n1369(net2283_c1,net2283);
INTERCONNECT GCLK_Pad_SplitCLK_0_1547(GCLK_Pad,net2284);
INTERCONNECT Split_HOLD_1667_DFFT_270__FPB_n1450(net2285_c1,net2285);
INTERCONNECT Split_HOLD_1668_DFFT_195__FPB_n1375(net2286_c1,net2286);
INTERCONNECT Split_HOLD_1669_DFFT_291__FPB_n1471(net2287_c1,net2287);
INTERCONNECT Split_HOLD_1670_DFFT_427__FPB_n1607(net2288_c1,net2288);
INTERCONNECT Split_HOLD_1671_DFFT_514__FPB_n1694(net2289_c1,net2289);
INTERCONNECT Split_HOLD_1672_DFFT_177__FPB_n1357(net2290_c1,net2290);
INTERCONNECT Split_HOLD_1673_DFFT_343__FPB_n1523(net2291_c1,net2291);
INTERCONNECT Split_HOLD_1674_DFFT_501__FPB_n1681(net2292_c1,net2292);
INTERCONNECT Split_HOLD_1675_DFFT_404__FPB_n1584(net2293_c1,net2293);
INTERCONNECT Split_HOLD_1676_DFFT_331__FPB_n1511(net2294_c1,net2294);
INTERCONNECT Split_HOLD_1677_DFFT_210__FPB_n1390(net2295_c1,net2295);
INTERCONNECT Split_HOLD_1678_DFFT_233__FPB_n1413(net2296_c1,net2296);
INTERCONNECT Split_HOLD_1679_DFFT_216__FPB_n1396(net2297_c1,net2297);
INTERCONNECT Split_HOLD_1680_DFFT_398__FPB_n1578(net2298_c1,net2298);
INTERCONNECT Split_HOLD_1681_DFFT_388__FPB_n1568(net2299_c1,net2299);
INTERCONNECT Split_HOLD_1682_DFFT_298__FPB_n1478(net2300_c1,net2300);
INTERCONNECT Split_HOLD_1683_DFFT_385__FPB_n1565(net2301_c1,net2301);
INTERCONNECT Split_HOLD_1684_DFFT_457__FPB_n1637(net2302_c1,net2302);
INTERCONNECT Split_HOLD_1685_AND2T_28_n28(net2303_c1,net2303);

endmodule
