
# Created      : Tue Apr 7 14:34:52 2020
# Platform     : Sahand.usc.edu
# User         : Ting-Ru Lin

VERSION 5.8 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.0100000 ;

CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS ON ;

SITE CoreSite
    CLASS CORE ;
    SIZE 1.000000 BY 160.000000 ; 
END CoreSite

LAYER M1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    WIDTH 4.400000 ;
    SPACING 5.600000 ;
    SPACING 0.090000 ENDOFLINE 0.090000 WITHIN 0.025000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.060000
      WIDTH  0.100000  0.100000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 10.00000 10.000000 ;
END M1

LAYER via1
    TYPE CUT ;
    SPACING 5.600000 ;
    WIDTH 4.400000 ;
END via1

LAYER M2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    WIDTH 4.400000 ;
    SPACING 5.600000 ;
    SPACING 0.090000 ENDOFLINE 0.090000 WITHIN 0.025000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.060000
      WIDTH  0.100000  0.100000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 10.00000 10.00000 ;
END M2

LAYER via2
    TYPE CUT ;
    SPACING 5.500000 ;
    WIDTH 4.500000 ;
END via2

LAYER M3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    WIDTH 4.400000 ;
    SPACING 5.600000 ;
    SPACING 0.090000 ENDOFLINE 0.090000 WITHIN 0.025000 ;
    SPACINGTABLE
    PARALLELRUNLENGTH
                       0.000000
      WIDTH  0.000000  0.060000
      WIDTH  0.100000  0.100000
      WIDTH  0.750000  0.250000
      WIDTH  1.500000  0.450000 ;
    PITCH 10.00000 10.000000 ;
END M3

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIA VIA12 DEFAULT 
    LAYER M1 ;
        RECT -2.20000 -2.20000 2.20000 2.20000 ;
    LAYER via1 ;
        RECT -2.20000 -2.20000 2.20000 2.20000 ;
    LAYER M2 ;
        RECT -2.20000 -2.20000 2.20000 2.20000 ;
END VIA12

VIA VIA23 DEFAULT 
    LAYER M2 ;
        RECT -2.20000 -2.20000 2.20000 2.20000 ;
    LAYER via2 ;
        RECT -2.20000 -2.20000 2.20000 2.20000 ;
    LAYER M3 ;
        RECT -2.20000 -2.20000 2.20000 2.20000 ;
END VIA23
MACRO PAD
    CLASS CORE ;
    FOREIGN PAD 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 100.000000 BY 120.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M1 ;
        RECT 27.000 12.500 73.000 107.500 ;
        LAYER M3 ;
        RECT 27.000 12.500 73.000 107.500 ;
	END
    END a
END PAD
MACRO LSmitll_AND2T
    CLASS CORE ;
    FOREIGN LSmitll_AND2T 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 100.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 12.800 17.200 17.200 ;
        END
    END a
    PIN b
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 82.800 52.800 87.200 57.200 ;
        END
    END b
    PIN q
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 82.800 12.800 87.200 17.200 ;
        END
    END q	
    PIN clk
         DIRECTION INOUT ;
         USE SIGNAL ;
         PORT
         LAYER M3 ;
         RECT 12.800 52.800 17.200 57.200 ;
         END
    END clk
END LSmitll_AND2T

MACRO LSmitll_XORT
    CLASS CORE ;
    FOREIGN LSmitll_XORT 0.000000 0.000000 ;	
    ORIGIN 0.000000 0.000000 ;
    SIZE 100.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 52.800 17.200 57.200 ;
        END
    END a
    PIN b
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 12.800 17.200 17.200 ;
        END
    END b
    PIN q
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 82.800 12.800 87.200 17.200 ;
        END
    END q	
    PIN clk
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 82.800 52.800 87.200 57.200 ;
        END
    END clk
END LSmitll_XORT

MACRO LSmitll_OR2T
    CLASS CORE ;
    FOREIGN LSmitll_XORT 0.000000 0.000000 ;	
    ORIGIN 0.000000 0.000000 ;
    SIZE 100.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 12.800 17.200 17.200 ;
        END
    END a
    PIN b
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 52.800 17.200 57.200 ;
        END
    END b
    PIN q
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 82.800 12.800 87.200 17.200 ;
        END
    END q	
    PIN clk
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 82.800 52.800 87.200 57.200 ;
        END
    END clk
END LSmitll_OR2T

MACRO LSmitll_NOTT
    CLASS CORE ;
    FOREIGN LSmitll_NOTT 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 100.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 52.800 17.200 57.200 ;
        END
    END a
    PIN q
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 82.800 12.800 87.200 17.200 ;
        END
    END q
    PIN clk
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 12.800 17.200 17.200 ;
        END
    END clk
END LSmitll_NOTT

MACRO LSmitll_DFFT
    CLASS CORE ;
    FOREIGN LSmitll_DFFT 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 80.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 12.800 17.200 17.200 ;
        END
    END a
    PIN q
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 62.800 12.800 67.200 17.200 ;
        END
    END q
    PIN clk
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 52.800 17.200 57.200 ;
        END
    END clk
END LSmitll_DFFT

MACRO LSmitll_NDROT
    CLASS CORE ;
    FOREIGN LSmitll_NDROT 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 120.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 52.800 17.200 57.200 ;
        END
    END a
	PIN b
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 12.800 17.200 17.200 ;
        END
    END b
    PIN q
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 102.800 12.800 107.200 17.200 ;
        END
    END q
    PIN clk
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 102.800 52.800 107.200 57.200 ;
        END
    END clk
END LSmitll_NDROT

MACRO LSmitll_SPLITT
    CLASS CORE ;
    FOREIGN LSmitll_SPLITT 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 50.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 52.800 17.200 57.200 ;
        END
    END a
    PIN q0
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 12.800 17.200 17.200 ;
        END
    END q0
    PIN q1
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 32.800 12.800 37.200 17.200 ;
        END
    END q1
END LSmitll_SPLITT

MACRO LSmitll_MERGET
    CLASS CORE ;
    FOREIGN LSmitll_MERGET 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 70.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ; 
    PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 12.800 17.200 17.200 ;
        END
    END a
    PIN b
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 12.800 52.800 17.200 57.200 ;
        END
    END b
    PIN q
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 62.800 12.800 67.200 17.200 ;
        END
    END q
END LSmitll_MERGET

MACRO LSmitll_JTLT
    CLASS CORE ;
    FOREIGN LSmitll_JTLT 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 40.000000 BY 70.000000 ;
    SYMMETRY X ;
    SITE CoreSite ;
	PIN a
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 2.800 52.800 7.200 57.200 ;
        END
    END a
    PIN q
        DIRECTION INOUT ;
        USE SIGNAL ;
        PORT
        LAYER M3 ;
        RECT 32.800 12.800 37.200 17.200 ;
        END
    END q
END LSmitll_JTLT

END LIBRARY

