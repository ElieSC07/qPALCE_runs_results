module TAP_route(
input GCLK_Pad,
input TMS_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output state_obs2_Pad,
output state_obs3_Pad);

wire TMS_Pad;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire TRST_Pad;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire state_obs0_Pad;
wire net461_c1;
wire state_obs1_Pad;
wire net462_c1;
wire state_obs2_Pad;
wire net463_c1;
wire state_obs3_Pad;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire net486_c1;
wire net486;
wire net487_c1;
wire net487;
wire net488_c1;
wire net488;
wire net489_c1;
wire net489;
wire net490_c1;
wire net490;
wire net491_c1;
wire net491;
wire net492_c1;
wire net492;
wire net493_c1;
wire net493;
wire net494_c1;
wire net494;
wire net495_c1;
wire net495;
wire net496_c1;
wire net496;
wire net497_c1;
wire net497;
wire net498_c1;
wire net498;
wire net499_c1;
wire net499;
wire net500_c1;
wire net500;
wire net501_c1;
wire net501;
wire net502_c1;
wire net502;
wire net503_c1;
wire net503;
wire net504_c1;
wire net504;
wire net505_c1;
wire net505;
wire net506_c1;
wire net506;
wire net507_c1;
wire net507;
wire net508_c1;
wire net508;
wire net509_c1;
wire net509;
wire net510_c1;
wire net510;
wire net511_c1;
wire net511;
wire net512_c1;
wire net512;
wire net513_c1;
wire net513;
wire net514_c1;
wire net514;
wire net515_c1;
wire net515;
wire net516_c1;
wire net516;
wire net517_c1;
wire net517;
wire net518_c1;
wire net518;
wire net519_c1;
wire net519;
wire net520_c1;
wire net520;
wire net521_c1;
wire net521;
wire net522_c1;
wire net522;
wire net523_c1;
wire net523;
wire net524_c1;
wire net524;
wire net525_c1;
wire net525;
wire net526_c1;
wire net526;
wire net527_c1;
wire net527;
wire net528_c1;
wire net528;
wire net529_c1;
wire net529;
wire net530_c1;
wire net530;
wire net531_c1;
wire net531;
wire net532_c1;
wire net532;
wire net533_c1;
wire net533;
wire net534_c1;
wire net534;
wire net535_c1;
wire net535;
wire net536_c1;
wire net536;
wire net537_c1;
wire net537;
wire net538_c1;
wire net538;
wire net539_c1;
wire net539;
wire net540_c1;
wire net540;
wire net541_c1;
wire net541;
wire net542_c1;
wire net542;
wire net543_c1;
wire net543;
wire net544_c1;
wire net544;
wire net545_c1;
wire net545;
wire net546_c1;
wire net546;
wire net547_c1;
wire net547;
wire net548_c1;
wire net548;
wire net549_c1;
wire net549;
wire net550_c1;
wire net550;
wire net551_c1;
wire net551;
wire net552_c1;
wire net552;
wire net553_c1;
wire net553;
wire net554_c1;
wire net554;
wire net555_c1;
wire net555;
wire net556_c1;
wire net556;
wire net557_c1;
wire net557;
wire net558_c1;
wire net558;
wire net559_c1;
wire net559;
wire net560_c1;
wire net560;
wire net561_c1;
wire net561;
wire net562_c1;
wire net562;
wire net563_c1;
wire net563;
wire net564_c1;
wire net564;
wire net565_c1;
wire net565;
wire net566_c1;
wire net566;
wire net567_c1;
wire net567;
wire net568_c1;
wire net568;
wire net569_c1;
wire net569;
wire net570_c1;
wire net570;
wire net571_c1;
wire net571;
wire net572_c1;
wire net572;
wire net573_c1;
wire net573;
wire net574_c1;
wire net574;
wire net575_c1;
wire net575;
wire net576_c1;
wire net576;
wire net577_c1;
wire net577;
wire net578_c1;
wire net578;
wire net579_c1;
wire net579;
wire net580_c1;
wire net580;
wire net581_c1;
wire net581;
wire net582_c1;
wire net582;
wire net583_c1;
wire net583;
wire net584_c1;
wire net584;
wire net585_c1;
wire net585;
wire net586_c1;
wire net586;
wire net587_c1;
wire net587;
wire net588_c1;
wire net588;
wire net589_c1;
wire net589;
wire net590_c1;
wire net590;
wire net591_c1;
wire net591;
wire net592_c1;
wire net592;
wire net593_c1;
wire net593;
wire net594_c1;
wire net594;
wire net595_c1;
wire net595;
wire net596_c1;
wire net596;
wire net597_c1;
wire net597;
wire net598_c1;
wire net598;
wire net599_c1;
wire net599;
wire net600_c1;
wire net600;
wire net601_c1;
wire net601;
wire net602_c1;
wire net602;
wire net603_c1;
wire net603;
wire net604_c1;
wire net604;
wire net605_c1;
wire net605;
wire net606_c1;
wire net606;
wire net607_c1;
wire net607;
wire net608_c1;
wire net608;
wire net609_c1;
wire net609;
wire net610_c1;
wire net610;
wire net611_c1;
wire net611;
wire net612_c1;
wire net612;
wire net613_c1;
wire net613;
wire net614_c1;
wire net614;
wire net615_c1;
wire net615;
wire net616_c1;
wire net616;
wire net617_c1;
wire net617;
wire net618_c1;
wire net618;
wire net619_c1;
wire net619;
wire net620_c1;
wire net620;
wire net621_c1;
wire net621;
wire net622_c1;
wire net622;
wire net623_c1;
wire net623;
wire net624_c1;
wire net624;
wire net625_c1;
wire net625;
wire net626_c1;
wire net626;
wire net627_c1;
wire net627;
wire net628_c1;
wire net628;
wire net629_c1;
wire net629;
wire net630_c1;
wire net630;
wire net631_c1;
wire net631;
wire net632_c1;
wire net632;
wire net633_c1;
wire net633;
wire net634_c1;
wire net634;
wire net635_c1;
wire net635;
wire net636_c1;
wire net636;
wire net637_c1;
wire net637;
wire net638_c1;
wire net638;
wire net639_c1;
wire net639;
wire net640_c1;
wire net640;
wire net641_c1;
wire net641;
wire net642_c1;
wire net642;
wire net643_c1;
wire net643;
wire net644_c1;
wire net644;
wire net645_c1;
wire net645;
wire net646_c1;
wire net646;
wire net647_c1;
wire net647;
wire net648_c1;
wire net648;
wire net649_c1;
wire net649;
wire net650_c1;
wire net650;
wire net651_c1;
wire net651;
wire net652_c1;
wire net652;
wire net653_c1;
wire net653;
wire net654_c1;
wire net654;
wire net655_c1;
wire net655;
wire net656_c1;
wire net656;
wire net657_c1;
wire net657;
wire net658_c1;
wire net658;
wire net659_c1;
wire net659;
wire net660_c1;
wire net660;
wire net661_c1;
wire net661;
wire net662_c1;
wire net662;
wire net663_c1;
wire net663;
wire net664_c1;
wire net664;
wire net665_c1;
wire net665;
wire net666_c1;
wire net666;
wire net667_c1;
wire net667;
wire net668_c1;
wire net668;
wire net669_c1;
wire net669;
wire net670_c1;
wire net670;
wire net671_c1;
wire net671;
wire net672_c1;
wire net672;
wire net673_c1;
wire net673;
wire net674_c1;
wire net674;
wire net675_c1;
wire net675;
wire net676_c1;
wire net676;
wire net677_c1;
wire net677;
wire net678_c1;
wire net678;
wire net679_c1;
wire net679;
wire net680_c1;
wire net680;
wire net681_c1;
wire net681;
wire net682_c1;
wire net682;
wire net683_c1;
wire net683;
wire net684_c1;
wire net684;
wire net685_c1;
wire net685;
wire net686_c1;
wire net686;
wire net687_c1;
wire net687;
wire net688_c1;
wire net688;
wire net689_c1;
wire net689;
wire net690_c1;
wire net690;
wire net691_c1;
wire net691;
wire net692_c1;
wire net692;
wire net693_c1;
wire net693;
wire net694_c1;
wire net694;
wire net695_c1;
wire net695;
wire net696_c1;
wire net696;
wire net697_c1;
wire net697;
wire net698_c1;
wire net698;
wire net699_c1;
wire net699;
wire net700_c1;
wire net700;
wire net701_c1;
wire net701;
wire net702_c1;
wire net702;
wire net703_c1;
wire net703;
wire net704_c1;
wire net704;
wire net705_c1;
wire net705;
wire net706_c1;
wire net706;
wire net707_c1;
wire net707;
wire net708_c1;
wire net708;
wire net709_c1;
wire net709;
wire net710_c1;
wire net710;
wire net711_c1;
wire net711;
wire net712_c1;
wire net712;
wire net713_c1;
wire net713;
wire net714_c1;
wire net714;
wire net715_c1;
wire net715;
wire net716_c1;
wire net716;
wire net717_c1;
wire net717;
wire net718_c1;
wire net718;
wire net719_c1;
wire net719;
wire net720_c1;
wire net720;
wire net721_c1;
wire net721;
wire net722_c1;
wire net722;
wire net723_c1;
wire net723;
wire net724_c1;
wire net724;
wire net725_c1;
wire net725;
wire net726_c1;
wire net726;
wire net727_c1;
wire net727;
wire net728_c1;
wire net728;
wire net729_c1;
wire net729;
wire net730_c1;
wire net730;
wire net731_c1;
wire net731;
wire net732_c1;
wire net732;
wire net733_c1;
wire net733;
wire net734_c1;
wire net734;
wire net735_c1;
wire net735;
wire net736_c1;
wire net736;
wire net737_c1;
wire net737;
wire net738_c1;
wire net738;
wire net739_c1;
wire net739;
wire net740_c1;
wire net740;
wire net741_c1;
wire net741;
wire net742_c1;
wire net742;
wire net743_c1;
wire net743;
wire net744_c1;
wire net744;
wire net745_c1;
wire net745;
wire net746_c1;
wire net746;
wire net747_c1;
wire net747;
wire net748_c1;
wire net748;
wire net749_c1;
wire net749;
wire net750_c1;
wire net750;
wire net751_c1;
wire net751;
wire net752_c1;
wire net752;
wire net753_c1;
wire net753;
wire net754_c1;
wire net754;
wire net755_c1;
wire net755;
wire net756_c1;
wire net756;
wire net757_c1;
wire net757;
wire net758_c1;
wire net758;
wire net759_c1;
wire net759;
wire net760_c1;
wire net760;
wire net761_c1;
wire net761;
wire net762_c1;
wire net762;
wire net763_c1;
wire net763;
wire net764_c1;
wire net764;
wire net765_c1;
wire net765;
wire net766_c1;
wire net766;
wire net767_c1;
wire net767;
wire net768_c1;
wire net768;
wire net769_c1;
wire net769;
wire net770_c1;
wire net770;
wire net771_c1;
wire net771;
wire net772_c1;
wire net772;
wire net773_c1;
wire net773;
wire net774_c1;
wire net774;
wire net775_c1;
wire net775;
wire net776_c1;
wire net776;
wire net777_c1;
wire net777;
wire net778_c1;
wire net778;
wire net779_c1;
wire net779;
wire net780_c1;
wire net780;
wire net781_c1;
wire net781;
wire net782_c1;
wire net782;
wire net783_c1;
wire net783;
wire net784_c1;
wire net784;
wire net785_c1;
wire net785;
wire net786_c1;
wire net786;
wire net787_c1;
wire net787;
wire net788_c1;
wire net788;
wire net789_c1;
wire net789;
wire net790_c1;
wire net790;
wire net791_c1;
wire net791;
wire net792_c1;
wire net792;
wire net793_c1;
wire net793;
wire net794_c1;
wire net794;
wire net795_c1;
wire net795;
wire net796_c1;
wire net796;
wire net797_c1;
wire net797;
wire net798_c1;
wire net798;
wire net799_c1;
wire net799;
wire net800_c1;
wire net800;
wire net801_c1;
wire net801;
wire net802_c1;
wire net802;
wire net803_c1;
wire net803;
wire net804_c1;
wire net804;
wire net805_c1;
wire net805;
wire net806_c1;
wire net806;
wire net807_c1;
wire net807;
wire net808_c1;
wire net808;
wire net809_c1;
wire net809;
wire net810_c1;
wire net810;
wire net811_c1;
wire net811;
wire net812_c1;
wire net812;
wire net813_c1;
wire net813;
wire net814_c1;
wire net814;
wire net815_c1;
wire net815;
wire net816_c1;
wire net816;
wire net817_c1;
wire net817;
wire net818_c1;
wire net818;
wire net819_c1;
wire net819;
wire net820_c1;
wire net820;
wire net821_c1;
wire net821;
wire net822_c1;
wire net822;
wire net823_c1;
wire net823;
wire net824_c1;
wire net824;
wire net825_c1;
wire net825;
wire net826_c1;
wire net826;
wire net827_c1;
wire net827;
wire net828_c1;
wire net828;
wire net829_c1;
wire net829;
wire net830_c1;
wire net830;
wire net831_c1;
wire net831;
wire net832_c1;
wire net832;
wire net833_c1;
wire net833;
wire net834_c1;
wire net834;
wire net835_c1;
wire net835;
wire net836_c1;
wire net836;
wire net837_c1;
wire net837;
wire net838_c1;
wire net838;
wire net839_c1;
wire net839;
wire net840_c1;
wire net840;
wire net841_c1;
wire net841;
wire net842_c1;
wire net842;
wire net843_c1;
wire net843;
wire net844_c1;
wire net844;
wire net845_c1;
wire net845;
wire net846_c1;
wire net846;
wire net847_c1;
wire net847;
wire net848_c1;
wire net848;
wire net849_c1;
wire net849;
wire net850_c1;
wire net850;
wire net851_c1;
wire net851;
wire net852_c1;
wire net852;
wire net853_c1;
wire net853;
wire net854_c1;
wire net854;
wire net855_c1;
wire net855;
wire net856_c1;
wire net856;
wire net857_c1;
wire net857;
wire net858_c1;
wire net858;
wire net859_c1;
wire net859;
wire net860_c1;
wire net860;
wire net861_c1;
wire net861;
wire net862_c1;
wire net862;
wire net863_c1;
wire net863;
wire net864_c1;
wire net864;
wire net865_c1;
wire net865;
wire net866_c1;
wire net866;
wire net867_c1;
wire net867;
wire net868_c1;
wire net868;
wire net869_c1;
wire net869;
wire net870_c1;
wire net870;
wire net871_c1;
wire net871;
wire net872_c1;
wire net872;
wire net873_c1;
wire net873;
wire net874_c1;
wire net874;
wire net875_c1;
wire net875;
wire net876_c1;
wire net876;
wire net877_c1;
wire net877;
wire net878_c1;
wire net878;
wire net879_c1;
wire net879;
wire net880_c1;
wire net880;
wire net881_c1;
wire net881;
wire net882_c1;
wire net882;
wire net883_c1;
wire net883;
wire net884_c1;
wire net884;
wire net885_c1;
wire net885;
wire net886_c1;
wire net886;
wire net887_c1;
wire net887;
wire net888_c1;
wire net888;
wire net889_c1;
wire net889;
wire net890_c1;
wire net890;
wire net891_c1;
wire net891;
wire net892_c1;
wire net892;
wire net893_c1;
wire net893;
wire net894_c1;
wire net894;
wire net895_c1;
wire net895;
wire net896_c1;
wire net896;
wire net897_c1;
wire net897;
wire net898_c1;
wire net898;
wire net899_c1;
wire net899;
wire net900_c1;
wire net900;
wire net901_c1;
wire net901;
wire net902_c1;
wire net902;
wire net903_c1;
wire net903;
wire net904_c1;
wire net904;
wire net905_c1;
wire net905;
wire net906_c1;
wire net906;
wire net907_c1;
wire net907;
wire net908_c1;
wire net908;
wire net909_c1;
wire net909;
wire net910_c1;
wire net910;
wire net911_c1;
wire net911;
wire net912_c1;
wire net912;
wire net913_c1;
wire net913;
wire net914_c1;
wire net914;
wire net915_c1;
wire net915;
wire net916_c1;
wire net916;
wire net917_c1;
wire net917;
wire net918_c1;
wire net918;
wire net919_c1;
wire net919;
wire net920_c1;
wire net920;
wire net921_c1;
wire net921;
wire net922_c1;
wire net922;
wire net923_c1;
wire net923;
wire net924_c1;
wire net924;
wire net925_c1;
wire net925;
wire net926_c1;
wire net926;
wire net927_c1;
wire net927;
wire net928_c1;
wire net928;
wire net929_c1;
wire net929;
wire net930_c1;
wire net930;
wire net931_c1;
wire net931;
wire net932_c1;
wire net932;
wire net933_c1;
wire net933;
wire net934_c1;
wire net934;
wire net935_c1;
wire net935;
wire net936_c1;
wire net936;
wire net937_c1;
wire net937;
wire net938_c1;
wire net938;
wire net939_c1;
wire net939;
wire net940_c1;
wire net940;
wire net941_c1;
wire net941;
wire net942_c1;
wire net942;
wire net943_c1;
wire net943;
wire net944_c1;
wire net944;
wire net945_c1;
wire net945;
wire net946_c1;
wire net946;
wire net947_c1;
wire net947;
wire net948_c1;
wire net948;
wire net949_c1;
wire net949;
wire net950_c1;
wire net950;
wire net951_c1;
wire net951;
wire net952_c1;
wire net952;
wire net953_c1;
wire net953;
wire net954_c1;
wire net954;
wire net955_c1;
wire net955;
wire net956_c1;
wire net956;
wire net957_c1;
wire net957;
wire net958_c1;
wire net958;
wire net959_c1;
wire net959;
wire net960_c1;
wire net960;
wire net961_c1;
wire net961;
wire net962_c1;
wire net962;
wire net963_c1;
wire net963;
wire net964_c1;
wire net964;
wire net965_c1;
wire net965;
wire net966_c1;
wire net966;
wire net967_c1;
wire net967;
wire net968_c1;
wire net968;
wire net969_c1;
wire net969;
wire net970_c1;
wire net970;
wire net971_c1;
wire net971;
wire GCLK_Pad;
wire net972;
wire net973_c1;
wire net973;
wire net974_c1;
wire net974;

DFFT DFFT_199__FPB_n592(net938,net433,net440_c1);
DFFT DFFT_241_state_obs0(net642,net384,net460_c1);
AND2T AND2T_101_n125(net876,net91,net358,net95_c1);
AND2T AND2T_110_n134(net870,net120,net395,net98_c1);
AND2T AND2T_102_n126(net924,net95,net362,net99_c1);
AND2T AND2T_103_n127(net888,net106,net366,net102_c1);
AND2T AND2T_122_n161(net622,net188,net281,net107_c1);
AND2T AND2T_114_n138(net690,net108,net388,net111_c1);
AND2T AND2T_107_n131(net948,net81,net381,net85_c1);
AND2T AND2T_108_n132(net902,net85,net102,net90_c1);
AND2T AND2T_109_n133(net768,net222,net389,net94_c1);
AND2T AND2T_125_n164(net674,net112,net403,net114_c1);
DFFT DFFT_254_state_obs2(net892,net425,net462_c1);
DFFT DFFT_248_state_obs1(net704,net376,net461_c1);
NOTT NOTT_8_n32(net748,net134,net2_c1);
NOTT NOTT_9_n33(net714,net316,net4_c1);
AND2T AND2T_10_n34(net684,net239,net408,net7_c1);
AND2T AND2T_20_n44(net762,net274,net390,net13_c1);
AND2T AND2T_12_n36(net816,net18,net359,net14_c1);
AND2T AND2T_21_n45(net778,net13,net398,net17_c1);
AND2T AND2T_13_n37(net817,net271,net363,net18_c1);
AND2T AND2T_30_n54(net564,net314,net174,net21_c1);
AND2T AND2T_14_n38(net800,net14,net369,net23_c1);
AND2T AND2T_31_n55(net752,net21,net290,net26_c1);
AND2T AND2T_16_n40(net826,net231,net375,net1_c1);
AND2T AND2T_40_n64(net784,net236,net159,net31_c1);
AND2T AND2T_24_n48(net776,net126,net254,net33_c1);
AND2T AND2T_17_n41(net889,net211,net297,net3_c1);
AND2T AND2T_41_n65(net827,net42,net415,net36_c1);
AND2T AND2T_25_n49(net764,net301,net251,net38_c1);
AND2T AND2T_26_n50(net566,net313,net416,net5_c1);
AND2T AND2T_50_n74(net496,net35,net414,net41_c1);
AND2T AND2T_34_n58(net698,net144,net368,net43_c1);
AND2T AND2T_19_n43(net567,net263,net383,net9_c1);
AND2T AND2T_51_n75(net608,net238,net422,net46_c1);
AND2T AND2T_43_n67(net574,net270,net423,net47_c1);
AND2T AND2T_35_n59(net576,net234,net199,net48_c1);
AND2T AND2T_36_n60(net502,net209,net243,net11_c1);
AND2T AND2T_28_n52(net620,net133,net250,net12_c1);
AND2T AND2T_60_n84(net769,net328,net405,net50_c1);
AND2T AND2T_52_n76(net670,net242,net128,net51_c1);
AND2T AND2T_44_n68(net588,net291,net129,net52_c1);
AND2T AND2T_29_n53(net668,net166,net252,net16_c1);
AND2T AND2T_53_n77(net691,net51,net46,net55_c1);
AND2T AND2T_45_n69(net550,net138,net228,net56_c1);
AND2T AND2T_38_n62(net794,net15,net397,net20_c1);
AND2T AND2T_54_n78(net682,net326,net437,net59_c1);
AND2T AND2T_39_n63(net777,net151,net406,net25_c1);
AND2T AND2T_55_n79(net824,net190,net220,net62_c1);
AND2T AND2T_56_n80(net832,net62,net442,net29_c1);
AND2T AND2T_64_n88(net512,net61,net421,net64_c1);
AND2T AND2T_66_n90(net520,net66,net441,net39_c1);
AND2T AND2T_58_n82(net590,net210,net447,net40_c1);
AND2T AND2T_74_n98(net575,net65,net449,net67_c1);
AND2T AND2T_67_n91(net763,net198,net450,net44_c1);
AND2T AND2T_59_n83(net770,net175,net396,net45_c1);
AND2T AND2T_68_n92(net582,net237,net266,net49_c1);
AND2T AND2T_69_n93(net771,net327,net412,net53_c1);
DFFT DFFT_259_state_obs3(net954,net399,net463_c1);
OR2T OR2T_22_n46(net754,net17,net23,net22_c1);
OR2T OR2T_23_n47(net551,net279,net407,net27_c1);
OR2T OR2T_32_n56(net765,net5,net424,net32_c1);
OR2T OR2T_33_n57(net746,net32,net22,net37_c1);
OR2T OR2T_42_n66(net825,net31,net325,net42_c1);
OR2T OR2T_37_n61(net490,net319,net374,net15_c1);
OR2T OR2T_61_n85(net596,net50,net40,net54_c1);
OR2T OR2T_46_n70(net565,net298,net431,net19_c1);
OR2T OR2T_70_n94(net583,net53,net49,net57_c1);
OR2T OR2T_62_n86(net597,net54,net34,net58_c1);
OR2T OR2T_47_n71(net801,net19,net36,net24_c1);
OR2T OR2T_71_n95(net580,net57,net44,net60_c1);
OR2T OR2T_63_n87(net518,net284,net413,net61_c1);
OR2T OR2T_48_n72(net755,net24,net20,net30_c1);
OR2T OR2T_72_n96(net532,net60,net39,net63_c1);
OR2T OR2T_57_n81(net594,net29,net59,net34_c1);
OR2T OR2T_49_n73(net747,net30,net37,net35_c1);
OR2T OR2T_73_n97(net534,net63,net58,net65_c1);
OR2T OR2T_65_n89(net514,net64,net215,net66_c1);
OR2T OR2T_75_n99(net846,net259,net453,net68_c1);
DFFT DFFT_130__PIPL_n181(net706,net465,net332_c1);
DFFT DFFT_131__PIPL_n182(net970,net113,net333_c1);
DFFT DFFT_132__PIPL_n183(net962,net89,net334_c1);
NOTT NOTT_11_n35(net840,net310,net10_c1);
NOTT NOTT_15_n39(net577,net267,net28_c1);
NOTT NOTT_18_n42(net814,net167,net6_c1);
NOTT NOTT_27_n51(net908,net191,net8_c1);
OR2T OR2T_100_n124(net862,net227,net324,net91_c1);
OR2T OR2T_111_n135(net858,net98,net94,net101_c1);
OR2T OR2T_112_n136(net864,net101,net404,net105_c1);
OR2T OR2T_104_n128(net886,net195,net218,net106_c1);
OR2T OR2T_113_n137(net877,net105,net99,net108_c1);
OR2T OR2T_105_n129(net964,net303,net287,net109_c1);
OR2T OR2T_106_n130(net955,net275,net373,net81_c1);
OR2T OR2T_116_n140(net900,net43,net394,net89_c1);
DFFT DFFT_117_state0_buf(net636,net143,net464_c1);
AND2T AND2T_80_n104(net830,net74,net80,net77_c1);
AND2T AND2T_81_n105(net920,net158,net448,net80_c1);
AND2T AND2T_90_n114(net595,net79,net285,net83_c1);
AND2T AND2T_91_n115(net688,net83,net458,net87_c1);
AND2T AND2T_84_n108(net612,net256,net452,net93_c1);
AND2T AND2T_77_n101(net934,net72,net457,net70_c1);
AND2T AND2T_85_n109(net614,net93,net454,net97_c1);
AND2T AND2T_86_n110(net628,net97,net456,net71_c1);
AND2T AND2T_78_n102(net940,net68,net440,net72_c1);
AND2T AND2T_79_n103(net831,net302,net300,net74_c1);
AND2T AND2T_95_n119(net941,net100,net367,net103_c1);
AND2T AND2T_88_n112(net720,net73,net307,net76_c1);
AND2T AND2T_98_n122(net901,net322,net241,net82_c1);
DFFT DFFT_129__PIPL_n180(net638,net464,net331_c1);
DFFT DFFT_200__FPB_n593(net925,net295,net444_c1);
DFFT DFFT_118_state1_buf(net699,net157,net465_c1);
DFFT DFFT_201__FPB_n594(net921,net444,net448_c1);
DFFT DFFT_210__FPB_n603(net796,net351,net354_c1);
DFFT DFFT_202__FPB_n595(net621,net160,net452_c1);
DFFT DFFT_211__FPB_n604(net797,net354,net357_c1);
DFFT DFFT_203__FPB_n596(net626,net88,net454_c1);
DFFT DFFT_140__FBL_n533(net926,net119,net338_c1);
DFFT DFFT_220__FPB_n613(net872,net78,net362_c1);
DFFT DFFT_212__FPB_n605(net810,net357,net361_c1);
DFFT DFFT_204__FPB_n597(net629,net84,net456_c1);
DFFT DFFT_141__FBL_n534(net675,net125,net339_c1);
DFFT DFFT_133__FBL_n526(net652,net317,net340_c1);
DFFT DFFT_221__FPB_n614(net700,net309,net366_c1);
DFFT DFFT_213__FPB_n606(net811,net361,net367_c1);
DFFT DFFT_205__FPB_n598(net715,net76,net458_c1);
DFFT DFFT_142__FBL_n535(net488,net213,net341_c1);
DFFT DFFT_134__FBL_n527(net535,net330,net342_c1);
DFFT DFFT_230__FPB_n623(net560,net365,net371_c1);
DFFT DFFT_222__FPB_n615(net650,net161,net373_c1);
DFFT DFFT_214__FPB_n607(net950,net194,net372_c1);
DFFT DFFT_150__FPB_n543(net838,net205,net375_c1);
DFFT DFFT_206__FPB_n599(net918,net77,net459_c1);
DFFT DFFT_143__FBL_n536(net528,net329,net343_c1);
DFFT DFFT_135__FBL_n528(net927,net226,net344_c1);
DFFT DFFT_207__FPB_n600(net932,net70,net348_c1);
DFFT DFFT_127__FPB_n178(net738,net156,net352_c1);
DFFT DFFT_231__FPB_n624(net561,net371,net378_c1);
DFFT DFFT_223__FPB_n616(net963,net974,net381_c1);
DFFT DFFT_215__FPB_n608(net949,net372,net382_c1);
DFFT DFFT_151__FPB_n544(net529,net315,net383_c1);
DFFT DFFT_144__FBL_n537(net951,net225,net345_c1);
DFFT DFFT_136__FBL_n529(net712,net233,net346_c1);
OR2T OR2T_82_n106(net651,net299,net132,net84_c1);
OR2T OR2T_83_n107(net627,net320,net149,net88_c1);
OR2T OR2T_76_n100(net919,net308,net455,net69_c1);
OR2T OR2T_92_n116(net676,net87,net71,net92_c1);
OR2T OR2T_93_n117(net878,net92,net459,net96_c1);
OR2T OR2T_94_n118(net935,net96,net348,net100_c1);
DFFT DFFT_208__FPB_n601(net749,net292,net349_c1);
DFFT DFFT_128__FPB_n179(net639,net268,net355_c1);
DFFT DFFT_240__FPB_n633(net643,net377,net384_c1);
DFFT DFFT_232__FPB_n625(net739,net378,net388_c1);
DFFT DFFT_224__FPB_n617(net685,net131,net389_c1);
DFFT DFFT_216__FPB_n609(net879,net186,net385_c1);
DFFT DFFT_160__FPB_n553(net808,net380,net387_c1);
DFFT DFFT_152__FPB_n545(net515,net249,net390_c1);
OR2T OR2T_87_n111(net658,net265,net246,net73_c1);
OR2T OR2T_96_n120(net833,net204,net196,net75_c1);
OR2T OR2T_97_n121(net871,net75,net219,net78_c1);
OR2T OR2T_89_n113(net591,net183,net269,net79_c1);
OR2T OR2T_99_n123(net689,net82,net382,net86_c1);
DFFT DFFT_137__FBL_n530(net503,net208,net335_c1);
DFFT DFFT_145__FBL_n538(net701,net230,net347_c1);
DFFT DFFT_217__FPB_n610(net903,net973,net350_c1);
DFFT DFFT_209__FPB_n602(net795,net349,net351_c1);
DFFT DFFT_233__FPB_n626(net894,net203,net394_c1);
DFFT DFFT_225__FPB_n618(net471,net221,net395_c1);
DFFT DFFT_161__FPB_n554(net802,net387,net397_c1);
DFFT DFFT_153__FPB_n546(net779,net293,net398_c1);
DFFT DFFT_138__FBL_n531(net521,net321,net336_c1);
DFFT DFFT_218__FPB_n611(net865,net350,net353_c1);
DFFT DFFT_250__FPB_n643(net906,net392,net400_c1);
DFFT DFFT_242__FPB_n635(net713,net332,net401_c1);
DFFT DFFT_234__FPB_n627(net677,net288,net403_c1);
DFFT DFFT_226__FPB_n619(net863,net90,net404_c1);
DFFT DFFT_170__FPB_n563(net484,net393,net402_c1);
DFFT DFFT_162__FPB_n555(net803,net171,net406_c1);
DFFT DFFT_154__FPB_n547(net504,net207,net407_c1);
DFFT DFFT_146__FPB_n539(net859,net305,net408_c1);
DFFT DFFT_139__FBL_n532(net526,net224,net337_c1);
DFFT DFFT_227__FPB_n620(net734,net185,net356_c1);
DFFT DFFT_219__FPB_n612(net887,net353,net358_c1);
DFFT DFFT_147__FPB_n540(net809,net121,net359_c1);
DFFT DFFT_251__FPB_n644(net907,net400,net409_c1);
DFFT DFFT_243__FPB_n636(net721,net401,net410_c1);
DFFT DFFT_235__FPB_n628(net644,net331,net411_c1);
DFFT DFFT_171__FPB_n564(net491,net402,net414_c1);
DFFT DFFT_163__FPB_n556(net844,net197,net415_c1);
DFFT DFFT_155__FPB_n548(net558,net182,net416_c1);
DFFT DFFT_228__FPB_n621(net735,net356,net360_c1);
DFFT DFFT_148__FPB_n541(net815,net276,net363_c1);
DFFT DFFT_252__FPB_n645(net895,net409,net417_c1);
DFFT DFFT_244__FPB_n637(net718,net410,net418_c1);
DFFT DFFT_236__FPB_n629(net656,net411,net419_c1);
DFFT DFFT_180__FPB_n573(net513,net142,net421_c1);
DFFT DFFT_172__FPB_n565(net609,net260,net422_c1);
DFFT DFFT_164__FPB_n557(net581,net272,net423_c1);
DFFT DFFT_156__FPB_n549(net740,net26,net424_c1);
DFFT DFFT_237__FPB_n630(net657,net419,net364_c1);
DFFT DFFT_229__FPB_n622(net470,net360,net365_c1);
DFFT DFFT_157__FPB_n550(net653,net214,net368_c1);
DFFT DFFT_149__FPB_n542(net753,net150,net369_c1);
DFFT DFFT_253__FPB_n646(net893,net417,net425_c1);
DFFT DFFT_245__FPB_n638(net719,net418,net426_c1);
DFFT DFFT_181__FPB_n574(net637,net136,net429_c1);
DFFT DFFT_173__FPB_n566(net613,net148,net430_c1);
DFFT DFFT_165__FPB_n558(net589,net56,net431_c1);
DFFT DFFT_238__FPB_n631(net659,net364,net370_c1);
DFFT DFFT_158__FPB_n551(net489,net11,net374_c1);
DFFT DFFT_246__FPB_n639(net707,net426,net432_c1);
DFFT DFFT_190__FPB_n583(net544,net428,net434_c1);
DFFT DFFT_182__FPB_n575(net469,net429,net435_c1);
DFFT DFFT_174__FPB_n567(net615,net430,net437_c1);
DFFT DFFT_166__FPB_n559(net498,net283,net436_c1);
SPLITT Split_300_n693(net306,net208_c1,net317_c1);
SPLITT Split_301_n694(net201,net213_c1,net321_c1);
SPLITT Split_310_n703(net111,net123_c1,net230_c1);
SPLITT Split_302_n695(net55,net217_c1,net324_c1);
SPLITT Split_311_n704(net123,net125_c1,net233_c1);
SPLITT Split_303_n696(net217,net219_c1,net326_c1);
SPLITT Split_312_n705(net115,net127_c1,net235_c1);
SPLITT Split_320_n713(net122,net128_c1,net236_c1);
SPLITT Split_304_n697(net45,net222_c1,net328_c1);
SPLITT Split_313_n706(net235,net133_c1,net239_c1);
SPLITT Split_321_n714(net107,net130_c1,net240_c1);
SPLITT Split_305_n698(net67,net223_c1,net329_c1);
SPLITT Split_314_n707(net127,net137_c1,net242_c1);
SPLITT Split_322_n715(net240,net138_c1,net243_c1);
SPLITT Split_330_n723(net117,net135_c1,net244_c1);
SPLITT Split_306_n699(net223,net224_c1,net330_c1);
SPLITT Split_307_n700(net103,net118_c1,net225_c1);
SPLITT Split_315_n708(net116,net140_c1,net248_c1);
SPLITT Split_323_n716(net130,net142_c1,net249_c1);
SPLITT Split_331_n724(net244,net144_c1,net250_c1);
SPLITT Split_308_n701(net118,net119_c1,net226_c1);
SPLITT Split_260_n653(net0,net147_c1,net253_c1);
SPLITT Split_316_n709(net248,net151_c1,net254_c1);
SPLITT Split_324_n717(net110,net146_c1,net255_c1);
SPLITT Split_332_n725(net135,net148_c1,net256_c1);
SPLITT Split_340_n733(net342,net145_c1,net257_c1);
SPLITT Split_309_n702(net86,net120_c1,net227_c1);
SPLITT Split_317_n710(net140,net121_c1,net228_c1);
SPLITT Split_261_n654(net253,net156_c1,net262_c1);
SPLITT Split_325_n718(net255,net159_c1,net263_c1);
SPLITT Split_333_n726(net352,net153_c1,net264_c1);
SPLITT Split_341_n734(net257,net157_c1,net265_c1);
SPLITT Split_318_n711(net104,net122_c1,net229_c1);
SPLITT Split_262_n655(net147,net161_c1,net268_c1);
SPLITT Split_270_n663(net154,net163_c1,net269_c1);
SPLITT Split_326_n719(net146,net165_c1,net270_c1);
SPLITT Split_334_n727(net264,net167_c1,net271_c1);
SPLITT Split_342_n735(net145,net160_c1,net272_c1);
SPLITT Split_350_n743(net338,net162_c1,net273_c1);
SPLITT Split_319_n712(net229,net126_c1,net231_c1);
SPLITT Split_327_n720(net114,net124_c1,net232_c1);
SPLITT Split_263_n656(net2,net169_c1,net277_c1);
SPLITT Split_271_n664(net28,net170_c1,net278_c1);
SPLITT Split_335_n728(net153,net174_c1,net279_c1);
SPLITT Split_343_n736(net344,net168_c1,net280_c1);
SPLITT Split_351_n744(net162,net172_c1,net281_c1);
SPLITT Split_328_n721(net232,net129_c1,net234_c1);
SPLITT Split_264_n657(net277,net180_c1,net283_c1);
SPLITT Split_272_n665(net170,net183_c1,net284_c1);
SPLITT Split_280_n673(net27,net182_c1,net285_c1);
SPLITT Split_336_n729(net355,net177_c1,net286_c1);
SPLITT Split_344_n737(net280,net181_c1,net287_c1);
SPLITT Split_352_n745(net339,net179_c1,net288_c1);
SPLITT Split_360_n753(net345,net176_c1,net289_c1);
SPLITT Split_329_n722(net124,net131_c1,net237_c1);
SPLITT Split_337_n730(net286,net132_c1,net238_c1);
SPLITT Split_265_n658(net169,net185_c1,net292_c1);
SPLITT Split_273_n666(net1,net187_c1,net293_c1);
SPLITT Split_281_n674(net33,net184_c1,net294_c1);
SPLITT Split_345_n738(net168,net186_c1,net295_c1);
SPLITT Split_353_n746(net179,net188_c1,net296_c1);
SPLITT Split_361_n754(net289,net191_c1,net297_c1);
DFFT DFFT_247__FPB_n640(net705,net432,net376_c1);
DFFT DFFT_239__FPB_n632(net645,net370,net377_c1);
DFFT DFFT_167__FPB_n560(net497,net436,net379_c1);
DFFT DFFT_159__FPB_n552(net741,net165,net380_c1);
SPLITT Split_338_n731(net177,net136_c1,net241_c1);
DFFT DFFT_255__FPB_n648(net956,net334,net438_c1);
DFFT DFFT_191__FPB_n584(net546,net434,net439_c1);
DFFT DFFT_183__FPB_n576(net533,net435,net441_c1);
DFFT DFFT_175__FPB_n568(net847,net312,net442_c1);
SPLITT Split_266_n659(net4,net195_c1,net299_c1);
SPLITT Split_274_n667(net187,net196_c1,net300_c1);
SPLITT Split_282_n675(net294,net199_c1,net301_c1);
SPLITT Split_290_n683(net178,net197_c1,net302_c1);
SPLITT Split_346_n739(net346,net194_c1,net303_c1);
SPLITT Split_354_n747(net341,net192_c1,net304_c1);
SPLITT Split_362_n755(net176,net193_c1,net305_c1);
SPLITT Split_267_n660(net7,net141_c1,net245_c1);
SPLITT Split_339_n732(net340,net143_c1,net246_c1);
SPLITT Split_347_n740(net336,net139_c1,net247_c1);
SPLITT Split_275_n668(net3,net203_c1,net307_c1);
SPLITT Split_283_n676(net184,net204_c1,net308_c1);
SPLITT Split_291_n684(net16,net202_c1,net309_c1);
SPLITT Split_355_n748(net304,net205_c1,net310_c1);
SPLITT Split_363_n756(net347,net200_c1,net311_c1);
SPLITT Split_268_n661(net141,net150_c1,net251_c1);
SPLITT Split_348_n741(net247,net149_c1,net252_c1);
SPLITT Split_276_n669(net6,net206_c1,net312_c1);
SPLITT Split_284_n677(net38,net210_c1,net313_c1);
SPLITT Split_292_n685(net202,net209_c1,net314_c1);
SPLITT Split_356_n749(net192,net207_c1,net315_c1);
SPLITT Split_364_n757(net311,net211_c1,net316_c1);
SPLITT Split_269_n662(net10,net154_c1,net258_c1);
SPLITT Split_277_n670(net206,net158_c1,net259_c1);
SPLITT Split_349_n742(net139,net155_c1,net260_c1);
SPLITT Split_357_n750(net343,net152_c1,net261_c1);
SPLITT Split_285_n678(net8,net212_c1,net318_c1);
SPLITT Split_293_n686(net48,net215_c1,net319_c1);
SPLITT Split_365_n758(net200,net214_c1,net320_c1);
SPLITT Split_278_n671(net9,net164_c1,net266_c1);
SPLITT Split_358_n751(net261,net166_c1,net267_c1);
SPLITT Split_286_n679(net318,net218_c1,net322_c1);
SPLITT Split_294_n687(net25,net216_c1,net323_c1);
SPLITT Split_279_n672(net164,net175_c1,net274_c1);
SPLITT Split_287_n680(net212,net173_c1,net275_c1);
SPLITT Split_359_n752(net152,net171_c1,net276_c1);
SPLITT Split_295_n688(net323,net220_c1,net325_c1);
SPLITT Split_288_n681(net12,net178_c1,net282_c1);
SPLITT Split_296_n689(net216,net221_c1,net327_c1);
SPLITT Split_289_n682(net282,net190_c1,net290_c1);
SPLITT Split_297_n690(net47,net189_c1,net291_c1);
SPLITT Split_298_n691(net52,net198_c1,net298_c1);
SPLITT Split_299_n692(net41,net201_c1,net306_c1);
NOTT NOTT_120_n159(net505,net335,net116_c1);
NOTT NOTT_121_n160(net527,net337,net104_c1);
NOTT NOTT_123_n162(net552,net262,net110_c1);
NOTT NOTT_115_n139(net968,net173,net113_c1);
NOTT NOTT_124_n163(net669,net172,net112_c1);
NOTT NOTT_126_n177(net623,net273,net117_c1);
NOTT NOTT_119_n158(net683,net296,net115_c1);
DFFT DFFT_168__FPB_n561(net485,net379,net386_c1);
DFFT DFFT_256__FPB_n649(net971,net438,net443_c1);
DFFT DFFT_192__FPB_n585(net559,net439,net445_c1);
DFFT DFFT_184__FPB_n577(net841,net163,net446_c1);
DFFT DFFT_176__FPB_n569(net553,net189,net447_c1);
DFFT DFFT_257__FPB_n650(net969,net443,net391_c1);
DFFT DFFT_249__FPB_n642(net909,net333,net392_c1);
DFFT DFFT_177__FPB_n570(net782,net278,net396_c1);
DFFT DFFT_169__FPB_n562(net468,net386,net393_c1);
DFFT DFFT_193__FPB_n586(net547,net445,net449_c1);
DFFT DFFT_185__FPB_n578(net839,net446,net450_c1);
DFFT DFFT_258__FPB_n651(net957,net391,net399_c1);
DFFT DFFT_178__FPB_n571(net783,net245,net405_c1);
DFFT DFFT_194__FPB_n587(net845,net258,net453_c1);
DFFT DFFT_186__FPB_n579(net873,net193,net451_c1);
DFFT DFFT_187__FPB_n580(net785,net451,net412_c1);
DFFT DFFT_179__FPB_n572(net519,net155,net413_c1);
DFFT DFFT_195__FPB_n588(net671,net137,net455_c1);
DFFT DFFT_188__FPB_n581(net499,net180,net420_c1);
DFFT DFFT_196__FPB_n589(net933,net69,net457_c1);
DFFT DFFT_197__FPB_n590(net965,net181,net427_c1);
DFFT DFFT_189__FPB_n582(net545,net420,net428_c1);
DFFT DFFT_198__FPB_n591(net939,net427,net433_c1);
SPLITT SplitCLK_4_253(net966,net971_c1,net970_c1);
SPLITT SplitCLK_4_254(net967,net969_c1,net968_c1);
SPLITT SplitCLK_4_255(net958,net967_c1,net966_c1);
SPLITT SplitCLK_4_256(net960,net965_c1,net964_c1);
SPLITT SplitCLK_0_257(net961,net962_c1,net963_c1);
SPLITT SplitCLK_0_258(net959,net961_c1,net960_c1);
SPLITT SplitCLK_4_259(net942,net958_c1,net959_c1);
SPLITT SplitCLK_4_260(net952,net956_c1,net957_c1);
SPLITT SplitCLK_4_261(net953,net954_c1,net955_c1);
SPLITT SplitCLK_6_262(net944,net952_c1,net953_c1);
SPLITT SplitCLK_4_263(net946,net951_c1,net950_c1);
SPLITT SplitCLK_4_264(net947,net948_c1,net949_c1);
SPLITT SplitCLK_4_265(net945,net947_c1,net946_c1);
SPLITT SplitCLK_2_266(net943,net945_c1,net944_c1);
SPLITT SplitCLK_6_267(net910,net942_c1,net943_c1);
SPLITT SplitCLK_4_268(net936,net941_c1,net940_c1);
SPLITT SplitCLK_0_269(net937,net938_c1,net939_c1);
SPLITT SplitCLK_0_270(net928,net937_c1,net936_c1);
SPLITT SplitCLK_4_271(net930,net934_c1,net935_c1);
SPLITT SplitCLK_4_272(net931,net932_c1,net933_c1);
SPLITT SplitCLK_6_273(net929,net930_c1,net931_c1);
SPLITT SplitCLK_4_274(net912,net929_c1,net928_c1);
SPLITT SplitCLK_4_275(net922,net927_c1,net926_c1);
SPLITT SplitCLK_4_276(net923,net924_c1,net925_c1);
SPLITT SplitCLK_6_277(net914,net922_c1,net923_c1);
SPLITT SplitCLK_4_278(net916,net920_c1,net921_c1);
SPLITT SplitCLK_4_279(net917,net919_c1,net918_c1);
SPLITT SplitCLK_4_280(net915,net917_c1,net916_c1);
SPLITT SplitCLK_2_281(net913,net915_c1,net914_c1);
SPLITT SplitCLK_4_282(net911,net913_c1,net912_c1);
SPLITT SplitCLK_0_283(net848,net910_c1,net911_c1);
SPLITT SplitCLK_4_284(net904,net908_c1,net909_c1);
SPLITT SplitCLK_4_285(net905,net907_c1,net906_c1);
SPLITT SplitCLK_6_286(net896,net904_c1,net905_c1);
SPLITT SplitCLK_4_287(net898,net903_c1,net902_c1);
SPLITT SplitCLK_4_288(net899,net901_c1,net900_c1);
SPLITT SplitCLK_2_289(net897,net898_c1,net899_c1);
SPLITT SplitCLK_0_290(net880,net896_c1,net897_c1);
SPLITT SplitCLK_4_291(net890,net894_c1,net895_c1);
SPLITT SplitCLK_4_292(net891,net892_c1,net893_c1);
SPLITT SplitCLK_6_293(net882,net890_c1,net891_c1);
SPLITT SplitCLK_4_294(net884,net889_c1,net888_c1);
SPLITT SplitCLK_4_295(net885,net886_c1,net887_c1);
SPLITT SplitCLK_4_296(net883,net885_c1,net884_c1);
SPLITT SplitCLK_2_297(net881,net883_c1,net882_c1);
SPLITT SplitCLK_6_298(net850,net880_c1,net881_c1);
SPLITT SplitCLK_4_299(net874,net879_c1,net878_c1);
SPLITT SplitCLK_4_300(net875,net876_c1,net877_c1);
SPLITT SplitCLK_4_301(net866,net875_c1,net874_c1);
SPLITT SplitCLK_4_302(net868,net873_c1,net872_c1);
SPLITT SplitCLK_4_303(net869,net871_c1,net870_c1);
SPLITT SplitCLK_4_304(net867,net869_c1,net868_c1);
SPLITT SplitCLK_0_305(net852,net866_c1,net867_c1);
SPLITT SplitCLK_4_306(net860,net865_c1,net864_c1);
SPLITT SplitCLK_4_307(net861,net863_c1,net862_c1);
SPLITT SplitCLK_2_308(net854,net860_c1,net861_c1);
SPLITT SplitCLK_4_309(net857,net859_c1,net858_c1);
SPLITT SplitCLK_4_310(net855,net856_c1,net857_c1);
SPLITT SplitCLK_2_311(net853,net855_c1,net854_c1);
SPLITT SplitCLK_4_312(net851,net853_c1,net852_c1);
SPLITT SplitCLK_2_313(net849,net851_c1,net850_c1);
SPLITT SplitCLK_6_314(net722,net848_c1,net849_c1);
SPLITT SplitCLK_4_315(net842,net846_c1,net847_c1);
SPLITT SplitCLK_4_316(net843,net845_c1,net844_c1);
SPLITT SplitCLK_6_317(net834,net842_c1,net843_c1);
SPLITT SplitCLK_4_318(net836,net841_c1,net840_c1);
SPLITT SplitCLK_4_319(net837,net838_c1,net839_c1);
SPLITT SplitCLK_4_320(net835,net837_c1,net836_c1);
SPLITT SplitCLK_0_321(net818,net834_c1,net835_c1);
SPLITT SplitCLK_4_322(net828,net833_c1,net832_c1);
SPLITT SplitCLK_4_323(net829,net831_c1,net830_c1);
SPLITT SplitCLK_2_324(net820,net828_c1,net829_c1);
SPLITT SplitCLK_4_325(net822,net826_c1,net827_c1);
SPLITT SplitCLK_4_326(net823,net825_c1,net824_c1);
SPLITT SplitCLK_4_327(net821,net823_c1,net822_c1);
SPLITT SplitCLK_2_328(net819,net821_c1,net820_c1);
SPLITT SplitCLK_6_329(net786,net818_c1,net819_c1);
SPLITT SplitCLK_4_330(net812,net816_c1,net817_c1);
SPLITT SplitCLK_0_331(net813,net814_c1,net815_c1);
SPLITT SplitCLK_6_332(net804,net812_c1,net813_c1);
SPLITT SplitCLK_4_333(net806,net810_c1,net811_c1);
SPLITT SplitCLK_4_334(net807,net808_c1,net809_c1);
SPLITT SplitCLK_4_335(net805,net807_c1,net806_c1);
SPLITT SplitCLK_4_336(net788,net804_c1,net805_c1);
SPLITT SplitCLK_4_337(net798,net803_c1,net802_c1);
SPLITT SplitCLK_4_338(net799,net801_c1,net800_c1);
SPLITT SplitCLK_6_339(net790,net798_c1,net799_c1);
SPLITT SplitCLK_4_340(net792,net796_c1,net797_c1);
SPLITT SplitCLK_2_341(net793,net795_c1,net794_c1);
SPLITT SplitCLK_4_342(net791,net793_c1,net792_c1);
SPLITT SplitCLK_2_343(net789,net791_c1,net790_c1);
SPLITT SplitCLK_4_344(net787,net789_c1,net788_c1);
SPLITT SplitCLK_0_345(net724,net786_c1,net787_c1);
SPLITT SplitCLK_4_346(net780,net785_c1,net784_c1);
SPLITT SplitCLK_4_347(net781,net782_c1,net783_c1);
SPLITT SplitCLK_2_348(net772,net781_c1,net780_c1);
SPLITT SplitCLK_4_349(net774,net778_c1,net779_c1);
SPLITT SplitCLK_4_350(net775,net777_c1,net776_c1);
SPLITT SplitCLK_4_351(net773,net775_c1,net774_c1);
SPLITT SplitCLK_6_352(net756,net773_c1,net772_c1);
SPLITT SplitCLK_4_353(net766,net771_c1,net770_c1);
SPLITT SplitCLK_4_354(net767,net768_c1,net769_c1);
SPLITT SplitCLK_6_355(net758,net766_c1,net767_c1);
SPLITT SplitCLK_4_356(net760,net765_c1,net764_c1);
SPLITT SplitCLK_4_357(net761,net762_c1,net763_c1);
SPLITT SplitCLK_2_358(net759,net760_c1,net761_c1);
SPLITT SplitCLK_6_359(net757,net758_c1,net759_c1);
SPLITT SplitCLK_6_360(net726,net756_c1,net757_c1);
SPLITT SplitCLK_4_361(net750,net755_c1,net754_c1);
SPLITT SplitCLK_0_362(net751,net752_c1,net753_c1);
SPLITT SplitCLK_0_363(net742,net751_c1,net750_c1);
SPLITT SplitCLK_4_364(net744,net749_c1,net748_c1);
SPLITT SplitCLK_4_365(net745,net746_c1,net747_c1);
SPLITT SplitCLK_4_366(net743,net745_c1,net744_c1);
SPLITT SplitCLK_4_367(net728,net742_c1,net743_c1);
SPLITT SplitCLK_4_368(net736,net741_c1,net740_c1);
SPLITT SplitCLK_4_369(net737,net739_c1,net738_c1);
SPLITT SplitCLK_4_370(net730,net737_c1,net736_c1);
SPLITT SplitCLK_4_371(net733,net735_c1,net734_c1);
SPLITT SplitCLK_4_372(net731,net732_c1,net733_c1);
SPLITT SplitCLK_6_373(net729,net730_c1,net731_c1);
SPLITT SplitCLK_4_374(net727,net729_c1,net728_c1);
SPLITT SplitCLK_4_375(net725,net726_c1,net727_c1);
SPLITT SplitCLK_4_376(net723,net725_c1,net724_c1);
SPLITT SplitCLK_0_377(net466,net722_c1,net723_c1);
SPLITT SplitCLK_4_378(net716,net720_c1,net721_c1);
SPLITT SplitCLK_4_379(net717,net719_c1,net718_c1);
SPLITT SplitCLK_6_380(net708,net716_c1,net717_c1);
SPLITT SplitCLK_4_381(net710,net715_c1,net714_c1);
SPLITT SplitCLK_4_382(net711,net713_c1,net712_c1);
SPLITT SplitCLK_4_383(net709,net711_c1,net710_c1);
SPLITT SplitCLK_0_384(net692,net708_c1,net709_c1);
SPLITT SplitCLK_4_385(net702,net706_c1,net707_c1);
SPLITT SplitCLK_4_386(net703,net704_c1,net705_c1);
SPLITT SplitCLK_6_387(net694,net702_c1,net703_c1);
SPLITT SplitCLK_4_388(net696,net700_c1,net701_c1);
SPLITT SplitCLK_4_389(net697,net698_c1,net699_c1);
SPLITT SplitCLK_2_390(net695,net696_c1,net697_c1);
SPLITT SplitCLK_2_391(net693,net695_c1,net694_c1);
SPLITT SplitCLK_6_392(net660,net692_c1,net693_c1);
SPLITT SplitCLK_4_393(net686,net690_c1,net691_c1);
SPLITT SplitCLK_4_394(net687,net688_c1,net689_c1);
SPLITT SplitCLK_2_395(net678,net686_c1,net687_c1);
SPLITT SplitCLK_4_396(net680,net685_c1,net684_c1);
SPLITT SplitCLK_4_397(net681,net682_c1,net683_c1);
SPLITT SplitCLK_4_398(net679,net681_c1,net680_c1);
SPLITT SplitCLK_0_399(net662,net678_c1,net679_c1);
SPLITT SplitCLK_4_400(net672,net676_c1,net677_c1);
SPLITT SplitCLK_4_401(net673,net675_c1,net674_c1);
SPLITT SplitCLK_4_402(net664,net673_c1,net672_c1);
SPLITT SplitCLK_4_403(net666,net671_c1,net670_c1);
SPLITT SplitCLK_4_404(net667,net668_c1,net669_c1);
SPLITT SplitCLK_4_405(net665,net667_c1,net666_c1);
SPLITT SplitCLK_6_406(net663,net664_c1,net665_c1);
SPLITT SplitCLK_4_407(net661,net663_c1,net662_c1);
SPLITT SplitCLK_0_408(net598,net660_c1,net661_c1);
SPLITT SplitCLK_4_409(net654,net658_c1,net659_c1);
SPLITT SplitCLK_4_410(net655,net656_c1,net657_c1);
SPLITT SplitCLK_6_411(net646,net654_c1,net655_c1);
SPLITT SplitCLK_4_412(net648,net652_c1,net653_c1);
SPLITT SplitCLK_4_413(net649,net650_c1,net651_c1);
SPLITT SplitCLK_2_414(net647,net648_c1,net649_c1);
SPLITT SplitCLK_6_415(net630,net647_c1,net646_c1);
SPLITT SplitCLK_4_416(net640,net644_c1,net645_c1);
SPLITT SplitCLK_0_417(net641,net642_c1,net643_c1);
SPLITT SplitCLK_6_418(net632,net640_c1,net641_c1);
SPLITT SplitCLK_4_419(net634,net639_c1,net638_c1);
SPLITT SplitCLK_4_420(net635,net636_c1,net637_c1);
SPLITT SplitCLK_6_421(net633,net634_c1,net635_c1);
SPLITT SplitCLK_6_422(net631,net632_c1,net633_c1);
SPLITT SplitCLK_6_423(net600,net630_c1,net631_c1);
SPLITT SplitCLK_4_424(net624,net629_c1,net628_c1);
SPLITT SplitCLK_4_425(net625,net626_c1,net627_c1);
SPLITT SplitCLK_6_426(net616,net624_c1,net625_c1);
SPLITT SplitCLK_4_427(net618,net623_c1,net622_c1);
SPLITT SplitCLK_4_428(net619,net620_c1,net621_c1);
SPLITT SplitCLK_4_429(net617,net619_c1,net618_c1);
SPLITT SplitCLK_0_430(net602,net616_c1,net617_c1);
SPLITT SplitCLK_4_431(net610,net614_c1,net615_c1);
SPLITT SplitCLK_0_432(net611,net612_c1,net613_c1);
SPLITT SplitCLK_0_433(net604,net611_c1,net610_c1);
SPLITT SplitCLK_4_434(net607,net608_c1,net609_c1);
SPLITT SplitCLK_2_435(net605,net606_c1,net607_c1);
SPLITT SplitCLK_4_436(net603,net605_c1,net604_c1);
SPLITT SplitCLK_4_437(net601,net603_c1,net602_c1);
SPLITT SplitCLK_6_438(net599,net600_c1,net601_c1);
SPLITT SplitCLK_6_439(net472,net598_c1,net599_c1);
SPLITT SplitCLK_4_440(net592,net597_c1,net596_c1);
SPLITT SplitCLK_4_441(net593,net594_c1,net595_c1);
SPLITT SplitCLK_6_442(net584,net592_c1,net593_c1);
SPLITT SplitCLK_4_443(net586,net591_c1,net590_c1);
SPLITT SplitCLK_4_444(net587,net588_c1,net589_c1);
SPLITT SplitCLK_4_445(net585,net587_c1,net586_c1);
SPLITT SplitCLK_4_446(net568,net585_c1,net584_c1);
SPLITT SplitCLK_4_447(net578,net583_c1,net582_c1);
SPLITT SplitCLK_4_448(net579,net581_c1,net580_c1);
SPLITT SplitCLK_6_449(net570,net578_c1,net579_c1);
SPLITT SplitCLK_4_450(net572,net576_c1,net577_c1);
SPLITT SplitCLK_4_451(net573,net574_c1,net575_c1);
SPLITT SplitCLK_6_452(net571,net572_c1,net573_c1);
SPLITT SplitCLK_6_453(net569,net570_c1,net571_c1);
SPLITT SplitCLK_2_454(net536,net568_c1,net569_c1);
SPLITT SplitCLK_4_455(net562,net567_c1,net566_c1);
SPLITT SplitCLK_4_456(net563,net565_c1,net564_c1);
SPLITT SplitCLK_6_457(net554,net562_c1,net563_c1);
SPLITT SplitCLK_4_458(net556,net561_c1,net560_c1);
SPLITT SplitCLK_4_459(net557,net559_c1,net558_c1);
SPLITT SplitCLK_4_460(net555,net557_c1,net556_c1);
SPLITT SplitCLK_0_461(net538,net554_c1,net555_c1);
SPLITT SplitCLK_4_462(net548,net553_c1,net552_c1);
SPLITT SplitCLK_0_463(net549,net550_c1,net551_c1);
SPLITT SplitCLK_4_464(net540,net549_c1,net548_c1);
SPLITT SplitCLK_4_465(net542,net547_c1,net546_c1);
SPLITT SplitCLK_4_466(net543,net545_c1,net544_c1);
SPLITT SplitCLK_4_467(net541,net543_c1,net542_c1);
SPLITT SplitCLK_6_468(net539,net540_c1,net541_c1);
SPLITT SplitCLK_4_469(net537,net539_c1,net538_c1);
SPLITT SplitCLK_4_470(net474,net536_c1,net537_c1);
SPLITT SplitCLK_4_471(net530,net535_c1,net534_c1);
SPLITT SplitCLK_4_472(net531,net533_c1,net532_c1);
SPLITT SplitCLK_6_473(net522,net530_c1,net531_c1);
SPLITT SplitCLK_4_474(net524,net529_c1,net528_c1);
SPLITT SplitCLK_0_475(net525,net526_c1,net527_c1);
SPLITT SplitCLK_0_476(net523,net525_c1,net524_c1);
SPLITT SplitCLK_0_477(net506,net522_c1,net523_c1);
SPLITT SplitCLK_4_478(net516,net521_c1,net520_c1);
SPLITT SplitCLK_4_479(net517,net518_c1,net519_c1);
SPLITT SplitCLK_6_480(net508,net516_c1,net517_c1);
SPLITT SplitCLK_4_481(net510,net514_c1,net515_c1);
SPLITT SplitCLK_4_482(net511,net512_c1,net513_c1);
SPLITT SplitCLK_4_483(net509,net511_c1,net510_c1);
SPLITT SplitCLK_2_484(net507,net509_c1,net508_c1);
SPLITT SplitCLK_6_485(net476,net506_c1,net507_c1);
SPLITT SplitCLK_4_486(net500,net504_c1,net505_c1);
SPLITT SplitCLK_4_487(net501,net502_c1,net503_c1);
SPLITT SplitCLK_4_488(net492,net501_c1,net500_c1);
SPLITT SplitCLK_4_489(net494,net498_c1,net499_c1);
SPLITT SplitCLK_2_490(net495,net497_c1,net496_c1);
SPLITT SplitCLK_4_491(net493,net495_c1,net494_c1);
SPLITT SplitCLK_4_492(net478,net493_c1,net492_c1);
SPLITT SplitCLK_4_493(net486,net490_c1,net491_c1);
SPLITT SplitCLK_4_494(net487,net488_c1,net489_c1);
SPLITT SplitCLK_2_495(net480,net486_c1,net487_c1);
SPLITT SplitCLK_4_496(net483,net484_c1,net485_c1);
SPLITT SplitCLK_2_497(net481,net482_c1,net483_c1);
SPLITT SplitCLK_2_498(net479,net481_c1,net480_c1);
SPLITT SplitCLK_4_499(net477,net479_c1,net478_c1);
SPLITT SplitCLK_2_500(net475,net477_c1,net476_c1);
SPLITT SplitCLK_4_501(net473,net475_c1,net474_c1);
SPLITT SplitCLK_2_502(net467,net473_c1,net472_c1);
wire dummy0;
SPLITT SplitCLK_2_503(net856,net471_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_2_504(net732,net470_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_505(net606,net469_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_506(net482,net468_c1,dummy3);
SPLITT SplitCLK_0_507(net972,net466_c1,net467_c1);
wire dummy4;
SPLITT Split_HOLD_621(net385,dummy4,net973_c1);
wire dummy5;
SPLITT Split_HOLD_622(net109,dummy5,net974_c1);
INTERCONNECT TMS_Pad_Split_260_n653(TMS_Pad,net0);
INTERCONNECT AND2T_16_n40_Split_273_n666(net1_c1,net1);
INTERCONNECT NOTT_8_n32_Split_263_n656(net2_c1,net2);
INTERCONNECT AND2T_17_n41_Split_275_n668(net3_c1,net3);
INTERCONNECT NOTT_9_n33_Split_266_n659(net4_c1,net4);
INTERCONNECT AND2T_26_n50_OR2T_32_n56(net5_c1,net5);
INTERCONNECT NOTT_18_n42_Split_276_n669(net6_c1,net6);
INTERCONNECT AND2T_10_n34_Split_267_n660(net7_c1,net7);
INTERCONNECT NOTT_27_n51_Split_285_n678(net8_c1,net8);
INTERCONNECT AND2T_19_n43_Split_278_n671(net9_c1,net9);
INTERCONNECT NOTT_11_n35_Split_269_n662(net10_c1,net10);
INTERCONNECT AND2T_36_n60_DFFT_158__FPB_n551(net11_c1,net11);
INTERCONNECT AND2T_28_n52_Split_288_n681(net12_c1,net12);
INTERCONNECT AND2T_20_n44_AND2T_21_n45(net13_c1,net13);
INTERCONNECT AND2T_12_n36_AND2T_14_n38(net14_c1,net14);
INTERCONNECT OR2T_37_n61_AND2T_38_n62(net15_c1,net15);
INTERCONNECT AND2T_29_n53_Split_291_n684(net16_c1,net16);
INTERCONNECT AND2T_21_n45_OR2T_22_n46(net17_c1,net17);
INTERCONNECT AND2T_13_n37_AND2T_12_n36(net18_c1,net18);
INTERCONNECT OR2T_46_n70_OR2T_47_n71(net19_c1,net19);
INTERCONNECT AND2T_38_n62_OR2T_48_n72(net20_c1,net20);
INTERCONNECT AND2T_30_n54_AND2T_31_n55(net21_c1,net21);
INTERCONNECT OR2T_22_n46_OR2T_33_n57(net22_c1,net22);
INTERCONNECT AND2T_14_n38_OR2T_22_n46(net23_c1,net23);
INTERCONNECT OR2T_47_n71_OR2T_48_n72(net24_c1,net24);
INTERCONNECT AND2T_39_n63_Split_294_n687(net25_c1,net25);
INTERCONNECT AND2T_31_n55_DFFT_156__FPB_n549(net26_c1,net26);
INTERCONNECT OR2T_23_n47_Split_280_n673(net27_c1,net27);
INTERCONNECT NOTT_15_n39_Split_271_n664(net28_c1,net28);
INTERCONNECT AND2T_56_n80_OR2T_57_n81(net29_c1,net29);
INTERCONNECT OR2T_48_n72_OR2T_49_n73(net30_c1,net30);
INTERCONNECT AND2T_40_n64_OR2T_42_n66(net31_c1,net31);
INTERCONNECT OR2T_32_n56_OR2T_33_n57(net32_c1,net32);
INTERCONNECT AND2T_24_n48_Split_281_n674(net33_c1,net33);
INTERCONNECT OR2T_57_n81_OR2T_62_n86(net34_c1,net34);
INTERCONNECT OR2T_49_n73_AND2T_50_n74(net35_c1,net35);
INTERCONNECT AND2T_41_n65_OR2T_47_n71(net36_c1,net36);
INTERCONNECT OR2T_33_n57_OR2T_49_n73(net37_c1,net37);
INTERCONNECT AND2T_25_n49_Split_284_n677(net38_c1,net38);
INTERCONNECT AND2T_66_n90_OR2T_72_n96(net39_c1,net39);
INTERCONNECT AND2T_58_n82_OR2T_61_n85(net40_c1,net40);
INTERCONNECT AND2T_50_n74_Split_299_n692(net41_c1,net41);
INTERCONNECT OR2T_42_n66_AND2T_41_n65(net42_c1,net42);
INTERCONNECT AND2T_34_n58_OR2T_116_n140(net43_c1,net43);
INTERCONNECT AND2T_67_n91_OR2T_71_n95(net44_c1,net44);
INTERCONNECT AND2T_59_n83_Split_304_n697(net45_c1,net45);
INTERCONNECT AND2T_51_n75_AND2T_53_n77(net46_c1,net46);
INTERCONNECT AND2T_43_n67_Split_297_n690(net47_c1,net47);
INTERCONNECT AND2T_35_n59_Split_293_n686(net48_c1,net48);
INTERCONNECT AND2T_68_n92_OR2T_70_n94(net49_c1,net49);
INTERCONNECT AND2T_60_n84_OR2T_61_n85(net50_c1,net50);
INTERCONNECT AND2T_52_n76_AND2T_53_n77(net51_c1,net51);
INTERCONNECT AND2T_44_n68_Split_298_n691(net52_c1,net52);
INTERCONNECT AND2T_69_n93_OR2T_70_n94(net53_c1,net53);
INTERCONNECT OR2T_61_n85_OR2T_62_n86(net54_c1,net54);
INTERCONNECT AND2T_53_n77_Split_302_n695(net55_c1,net55);
INTERCONNECT AND2T_45_n69_DFFT_165__FPB_n558(net56_c1,net56);
INTERCONNECT OR2T_70_n94_OR2T_71_n95(net57_c1,net57);
INTERCONNECT OR2T_62_n86_OR2T_73_n97(net58_c1,net58);
INTERCONNECT AND2T_54_n78_OR2T_57_n81(net59_c1,net59);
INTERCONNECT OR2T_71_n95_OR2T_72_n96(net60_c1,net60);
INTERCONNECT OR2T_63_n87_AND2T_64_n88(net61_c1,net61);
INTERCONNECT AND2T_55_n79_AND2T_56_n80(net62_c1,net62);
INTERCONNECT OR2T_72_n96_OR2T_73_n97(net63_c1,net63);
INTERCONNECT AND2T_64_n88_OR2T_65_n89(net64_c1,net64);
INTERCONNECT OR2T_73_n97_AND2T_74_n98(net65_c1,net65);
INTERCONNECT OR2T_65_n89_AND2T_66_n90(net66_c1,net66);
INTERCONNECT AND2T_74_n98_Split_305_n698(net67_c1,net67);
INTERCONNECT OR2T_75_n99_AND2T_78_n102(net68_c1,net68);
INTERCONNECT OR2T_76_n100_DFFT_196__FPB_n589(net69_c1,net69);
INTERCONNECT AND2T_77_n101_DFFT_207__FPB_n600(net70_c1,net70);
INTERCONNECT AND2T_86_n110_OR2T_92_n116(net71_c1,net71);
INTERCONNECT AND2T_78_n102_AND2T_77_n101(net72_c1,net72);
INTERCONNECT OR2T_87_n111_AND2T_88_n112(net73_c1,net73);
INTERCONNECT AND2T_79_n103_AND2T_80_n104(net74_c1,net74);
INTERCONNECT OR2T_96_n120_OR2T_97_n121(net75_c1,net75);
INTERCONNECT AND2T_88_n112_DFFT_205__FPB_n598(net76_c1,net76);
INTERCONNECT AND2T_80_n104_DFFT_206__FPB_n599(net77_c1,net77);
INTERCONNECT OR2T_97_n121_DFFT_220__FPB_n613(net78_c1,net78);
INTERCONNECT OR2T_89_n113_AND2T_90_n114(net79_c1,net79);
INTERCONNECT AND2T_81_n105_AND2T_80_n104(net80_c1,net80);
INTERCONNECT OR2T_106_n130_AND2T_107_n131(net81_c1,net81);
INTERCONNECT AND2T_98_n122_OR2T_99_n123(net82_c1,net82);
INTERCONNECT AND2T_90_n114_AND2T_91_n115(net83_c1,net83);
INTERCONNECT OR2T_82_n106_DFFT_204__FPB_n597(net84_c1,net84);
INTERCONNECT AND2T_107_n131_AND2T_108_n132(net85_c1,net85);
INTERCONNECT OR2T_99_n123_Split_309_n702(net86_c1,net86);
INTERCONNECT AND2T_91_n115_OR2T_92_n116(net87_c1,net87);
INTERCONNECT OR2T_83_n107_DFFT_203__FPB_n596(net88_c1,net88);
INTERCONNECT OR2T_116_n140_DFFT_132__PIPL_n183(net89_c1,net89);
INTERCONNECT AND2T_108_n132_DFFT_226__FPB_n619(net90_c1,net90);
INTERCONNECT OR2T_100_n124_AND2T_101_n125(net91_c1,net91);
INTERCONNECT OR2T_92_n116_OR2T_93_n117(net92_c1,net92);
INTERCONNECT AND2T_84_n108_AND2T_85_n109(net93_c1,net93);
INTERCONNECT AND2T_109_n133_OR2T_111_n135(net94_c1,net94);
INTERCONNECT AND2T_101_n125_AND2T_102_n126(net95_c1,net95);
INTERCONNECT OR2T_93_n117_OR2T_94_n118(net96_c1,net96);
INTERCONNECT AND2T_85_n109_AND2T_86_n110(net97_c1,net97);
INTERCONNECT AND2T_110_n134_OR2T_111_n135(net98_c1,net98);
INTERCONNECT AND2T_102_n126_OR2T_113_n137(net99_c1,net99);
INTERCONNECT OR2T_94_n118_AND2T_95_n119(net100_c1,net100);
INTERCONNECT OR2T_111_n135_OR2T_112_n136(net101_c1,net101);
INTERCONNECT AND2T_103_n127_AND2T_108_n132(net102_c1,net102);
INTERCONNECT AND2T_95_n119_Split_307_n700(net103_c1,net103);
INTERCONNECT NOTT_121_n160_Split_318_n711(net104_c1,net104);
INTERCONNECT OR2T_112_n136_OR2T_113_n137(net105_c1,net105);
INTERCONNECT OR2T_104_n128_AND2T_103_n127(net106_c1,net106);
INTERCONNECT AND2T_122_n161_Split_321_n714(net107_c1,net107);
INTERCONNECT OR2T_113_n137_AND2T_114_n138(net108_c1,net108);
INTERCONNECT OR2T_105_n129_Split_HOLD_622(net109_c1,net109);
INTERCONNECT NOTT_123_n162_Split_324_n717(net110_c1,net110);
INTERCONNECT AND2T_114_n138_Split_310_n703(net111_c1,net111);
INTERCONNECT NOTT_124_n163_AND2T_125_n164(net112_c1,net112);
INTERCONNECT NOTT_115_n139_DFFT_131__PIPL_n182(net113_c1,net113);
INTERCONNECT AND2T_125_n164_Split_327_n720(net114_c1,net114);
INTERCONNECT NOTT_119_n158_Split_312_n705(net115_c1,net115);
INTERCONNECT NOTT_120_n159_Split_315_n708(net116_c1,net116);
INTERCONNECT NOTT_126_n177_Split_330_n723(net117_c1,net117);
INTERCONNECT Split_307_n700_Split_308_n701(net118_c1,net118);
INTERCONNECT Split_308_n701_DFFT_140__FBL_n533(net119_c1,net119);
INTERCONNECT Split_309_n702_AND2T_110_n134(net120_c1,net120);
INTERCONNECT Split_317_n710_DFFT_147__FPB_n540(net121_c1,net121);
INTERCONNECT Split_318_n711_Split_320_n713(net122_c1,net122);
INTERCONNECT Split_310_n703_Split_311_n704(net123_c1,net123);
INTERCONNECT Split_327_n720_Split_329_n722(net124_c1,net124);
INTERCONNECT Split_311_n704_DFFT_141__FBL_n534(net125_c1,net125);
INTERCONNECT Split_319_n712_AND2T_24_n48(net126_c1,net126);
INTERCONNECT Split_312_n705_Split_314_n707(net127_c1,net127);
INTERCONNECT Split_320_n713_AND2T_52_n76(net128_c1,net128);
INTERCONNECT Split_328_n721_AND2T_44_n68(net129_c1,net129);
INTERCONNECT Split_321_n714_Split_323_n716(net130_c1,net130);
INTERCONNECT Split_329_n722_DFFT_224__FPB_n617(net131_c1,net131);
INTERCONNECT Split_337_n730_OR2T_82_n106(net132_c1,net132);
INTERCONNECT Split_313_n706_AND2T_28_n52(net133_c1,net133);
INTERCONNECT TRST_Pad_NOTT_8_n32(TRST_Pad,net134);
INTERCONNECT Split_330_n723_Split_332_n725(net135_c1,net135);
INTERCONNECT Split_338_n731_DFFT_181__FPB_n574(net136_c1,net136);
INTERCONNECT Split_314_n707_DFFT_195__FPB_n588(net137_c1,net137);
INTERCONNECT Split_322_n715_AND2T_45_n69(net138_c1,net138);
INTERCONNECT Split_347_n740_Split_349_n742(net139_c1,net139);
INTERCONNECT Split_315_n708_Split_317_n710(net140_c1,net140);
INTERCONNECT Split_267_n660_Split_268_n661(net141_c1,net141);
INTERCONNECT Split_323_n716_DFFT_180__FPB_n573(net142_c1,net142);
INTERCONNECT Split_339_n732_DFFT_117_state0_buf(net143_c1,net143);
INTERCONNECT Split_331_n724_AND2T_34_n58(net144_c1,net144);
INTERCONNECT Split_340_n733_Split_342_n735(net145_c1,net145);
INTERCONNECT Split_324_n717_Split_326_n719(net146_c1,net146);
INTERCONNECT Split_260_n653_Split_262_n655(net147_c1,net147);
INTERCONNECT Split_332_n725_DFFT_173__FPB_n566(net148_c1,net148);
INTERCONNECT Split_348_n741_OR2T_83_n107(net149_c1,net149);
INTERCONNECT Split_268_n661_DFFT_149__FPB_n542(net150_c1,net150);
INTERCONNECT Split_316_n709_AND2T_39_n63(net151_c1,net151);
INTERCONNECT Split_357_n750_Split_359_n752(net152_c1,net152);
INTERCONNECT Split_333_n726_Split_335_n728(net153_c1,net153);
INTERCONNECT Split_269_n662_Split_270_n663(net154_c1,net154);
INTERCONNECT Split_349_n742_DFFT_179__FPB_n572(net155_c1,net155);
INTERCONNECT Split_261_n654_DFFT_127__FPB_n178(net156_c1,net156);
INTERCONNECT Split_341_n734_DFFT_118_state1_buf(net157_c1,net157);
INTERCONNECT Split_277_n670_AND2T_81_n105(net158_c1,net158);
INTERCONNECT Split_325_n718_AND2T_40_n64(net159_c1,net159);
INTERCONNECT Split_342_n735_DFFT_202__FPB_n595(net160_c1,net160);
INTERCONNECT Split_262_n655_DFFT_222__FPB_n615(net161_c1,net161);
INTERCONNECT Split_350_n743_Split_351_n744(net162_c1,net162);
INTERCONNECT Split_270_n663_DFFT_184__FPB_n577(net163_c1,net163);
INTERCONNECT Split_278_n671_Split_279_n672(net164_c1,net164);
INTERCONNECT Split_326_n719_DFFT_159__FPB_n552(net165_c1,net165);
INTERCONNECT Split_358_n751_AND2T_29_n53(net166_c1,net166);
INTERCONNECT Split_334_n727_NOTT_18_n42(net167_c1,net167);
INTERCONNECT Split_343_n736_Split_345_n738(net168_c1,net168);
INTERCONNECT Split_263_n656_Split_265_n658(net169_c1,net169);
INTERCONNECT Split_271_n664_Split_272_n665(net170_c1,net170);
INTERCONNECT Split_359_n752_DFFT_162__FPB_n555(net171_c1,net171);
INTERCONNECT Split_351_n744_NOTT_124_n163(net172_c1,net172);
INTERCONNECT Split_287_n680_NOTT_115_n139(net173_c1,net173);
INTERCONNECT Split_335_n728_AND2T_30_n54(net174_c1,net174);
INTERCONNECT Split_279_n672_AND2T_59_n83(net175_c1,net175);
INTERCONNECT Split_360_n753_Split_362_n755(net176_c1,net176);
INTERCONNECT Split_336_n729_Split_338_n731(net177_c1,net177);
INTERCONNECT Split_288_n681_Split_290_n683(net178_c1,net178);
INTERCONNECT Split_352_n745_Split_353_n746(net179_c1,net179);
INTERCONNECT Split_264_n657_DFFT_188__FPB_n581(net180_c1,net180);
INTERCONNECT Split_344_n737_DFFT_197__FPB_n590(net181_c1,net181);
INTERCONNECT Split_280_n673_DFFT_155__FPB_n548(net182_c1,net182);
INTERCONNECT Split_272_n665_OR2T_89_n113(net183_c1,net183);
INTERCONNECT Split_281_n674_Split_283_n676(net184_c1,net184);
INTERCONNECT Split_265_n658_DFFT_227__FPB_n620(net185_c1,net185);
INTERCONNECT Split_345_n738_DFFT_216__FPB_n609(net186_c1,net186);
INTERCONNECT Split_273_n666_Split_274_n667(net187_c1,net187);
INTERCONNECT Split_353_n746_AND2T_122_n161(net188_c1,net188);
INTERCONNECT Split_297_n690_DFFT_176__FPB_n569(net189_c1,net189);
INTERCONNECT Split_289_n682_AND2T_55_n79(net190_c1,net190);
INTERCONNECT Split_361_n754_NOTT_27_n51(net191_c1,net191);
INTERCONNECT Split_354_n747_Split_356_n749(net192_c1,net192);
INTERCONNECT Split_362_n755_DFFT_186__FPB_n579(net193_c1,net193);
INTERCONNECT Split_346_n739_DFFT_214__FPB_n607(net194_c1,net194);
INTERCONNECT Split_266_n659_OR2T_104_n128(net195_c1,net195);
INTERCONNECT Split_274_n667_OR2T_96_n120(net196_c1,net196);
INTERCONNECT Split_290_n683_DFFT_163__FPB_n556(net197_c1,net197);
INTERCONNECT Split_298_n691_AND2T_67_n91(net198_c1,net198);
INTERCONNECT Split_282_n675_AND2T_35_n59(net199_c1,net199);
INTERCONNECT Split_363_n756_Split_365_n758(net200_c1,net200);
INTERCONNECT Split_299_n692_Split_301_n694(net201_c1,net201);
INTERCONNECT Split_291_n684_Split_292_n685(net202_c1,net202);
INTERCONNECT Split_275_n668_DFFT_233__FPB_n626(net203_c1,net203);
INTERCONNECT Split_283_n676_OR2T_96_n120(net204_c1,net204);
INTERCONNECT Split_355_n748_DFFT_150__FPB_n543(net205_c1,net205);
INTERCONNECT Split_276_n669_Split_277_n670(net206_c1,net206);
INTERCONNECT Split_356_n749_DFFT_154__FPB_n547(net207_c1,net207);
INTERCONNECT Split_300_n693_DFFT_137__FBL_n530(net208_c1,net208);
INTERCONNECT Split_292_n685_AND2T_36_n60(net209_c1,net209);
INTERCONNECT Split_284_n677_AND2T_58_n82(net210_c1,net210);
INTERCONNECT Split_364_n757_AND2T_17_n41(net211_c1,net211);
INTERCONNECT Split_285_n678_Split_287_n680(net212_c1,net212);
INTERCONNECT Split_301_n694_DFFT_142__FBL_n535(net213_c1,net213);
INTERCONNECT Split_365_n758_DFFT_157__FPB_n550(net214_c1,net214);
INTERCONNECT Split_293_n686_OR2T_65_n89(net215_c1,net215);
INTERCONNECT Split_294_n687_Split_296_n689(net216_c1,net216);
INTERCONNECT Split_302_n695_Split_303_n696(net217_c1,net217);
INTERCONNECT Split_286_n679_OR2T_104_n128(net218_c1,net218);
INTERCONNECT Split_303_n696_OR2T_97_n121(net219_c1,net219);
INTERCONNECT Split_295_n688_AND2T_55_n79(net220_c1,net220);
INTERCONNECT Split_296_n689_DFFT_225__FPB_n618(net221_c1,net221);
INTERCONNECT Split_304_n697_AND2T_109_n133(net222_c1,net222);
INTERCONNECT Split_305_n698_Split_306_n699(net223_c1,net223);
INTERCONNECT Split_306_n699_DFFT_139__FBL_n532(net224_c1,net224);
INTERCONNECT Split_307_n700_DFFT_144__FBL_n537(net225_c1,net225);
INTERCONNECT Split_308_n701_DFFT_135__FBL_n528(net226_c1,net226);
INTERCONNECT Split_309_n702_OR2T_100_n124(net227_c1,net227);
INTERCONNECT Split_317_n710_AND2T_45_n69(net228_c1,net228);
INTERCONNECT Split_318_n711_Split_319_n712(net229_c1,net229);
INTERCONNECT Split_310_n703_DFFT_145__FBL_n538(net230_c1,net230);
INTERCONNECT Split_319_n712_AND2T_16_n40(net231_c1,net231);
INTERCONNECT Split_327_n720_Split_328_n721(net232_c1,net232);
INTERCONNECT Split_311_n704_DFFT_136__FBL_n529(net233_c1,net233);
INTERCONNECT Split_328_n721_AND2T_35_n59(net234_c1,net234);
INTERCONNECT Split_312_n705_Split_313_n706(net235_c1,net235);
INTERCONNECT Split_320_n713_AND2T_40_n64(net236_c1,net236);
INTERCONNECT Split_329_n722_AND2T_68_n92(net237_c1,net237);
INTERCONNECT Split_337_n730_AND2T_51_n75(net238_c1,net238);
INTERCONNECT Split_313_n706_AND2T_10_n34(net239_c1,net239);
INTERCONNECT Split_321_n714_Split_322_n715(net240_c1,net240);
INTERCONNECT Split_338_n731_AND2T_98_n122(net241_c1,net241);
INTERCONNECT Split_314_n707_AND2T_52_n76(net242_c1,net242);
INTERCONNECT Split_322_n715_AND2T_36_n60(net243_c1,net243);
INTERCONNECT Split_330_n723_Split_331_n724(net244_c1,net244);
INTERCONNECT Split_267_n660_DFFT_178__FPB_n571(net245_c1,net245);
INTERCONNECT Split_339_n732_OR2T_87_n111(net246_c1,net246);
INTERCONNECT Split_347_n740_Split_348_n741(net247_c1,net247);
INTERCONNECT Split_315_n708_Split_316_n709(net248_c1,net248);
INTERCONNECT Split_323_n716_DFFT_152__FPB_n545(net249_c1,net249);
INTERCONNECT Split_331_n724_AND2T_28_n52(net250_c1,net250);
INTERCONNECT Split_268_n661_AND2T_25_n49(net251_c1,net251);
INTERCONNECT Split_348_n741_AND2T_29_n53(net252_c1,net252);
INTERCONNECT Split_260_n653_Split_261_n654(net253_c1,net253);
INTERCONNECT Split_316_n709_AND2T_24_n48(net254_c1,net254);
INTERCONNECT Split_324_n717_Split_325_n718(net255_c1,net255);
INTERCONNECT Split_332_n725_AND2T_84_n108(net256_c1,net256);
INTERCONNECT Split_340_n733_Split_341_n734(net257_c1,net257);
INTERCONNECT Split_269_n662_DFFT_194__FPB_n587(net258_c1,net258);
INTERCONNECT Split_277_n670_OR2T_75_n99(net259_c1,net259);
INTERCONNECT Split_349_n742_DFFT_172__FPB_n565(net260_c1,net260);
INTERCONNECT Split_357_n750_Split_358_n751(net261_c1,net261);
INTERCONNECT Split_261_n654_NOTT_123_n162(net262_c1,net262);
INTERCONNECT Split_325_n718_AND2T_19_n43(net263_c1,net263);
INTERCONNECT Split_333_n726_Split_334_n727(net264_c1,net264);
INTERCONNECT Split_341_n734_OR2T_87_n111(net265_c1,net265);
INTERCONNECT Split_278_n671_AND2T_68_n92(net266_c1,net266);
INTERCONNECT Split_358_n751_NOTT_15_n39(net267_c1,net267);
INTERCONNECT Split_262_n655_DFFT_128__FPB_n179(net268_c1,net268);
INTERCONNECT Split_270_n663_OR2T_89_n113(net269_c1,net269);
INTERCONNECT Split_326_n719_AND2T_43_n67(net270_c1,net270);
INTERCONNECT Split_334_n727_AND2T_13_n37(net271_c1,net271);
INTERCONNECT Split_342_n735_DFFT_164__FPB_n557(net272_c1,net272);
INTERCONNECT Split_350_n743_NOTT_126_n177(net273_c1,net273);
INTERCONNECT Split_279_n672_AND2T_20_n44(net274_c1,net274);
INTERCONNECT Split_287_n680_OR2T_106_n130(net275_c1,net275);
INTERCONNECT Split_359_n752_DFFT_148__FPB_n541(net276_c1,net276);
INTERCONNECT Split_263_n656_Split_264_n657(net277_c1,net277);
INTERCONNECT Split_271_n664_DFFT_177__FPB_n570(net278_c1,net278);
INTERCONNECT Split_335_n728_OR2T_23_n47(net279_c1,net279);
INTERCONNECT Split_343_n736_Split_344_n737(net280_c1,net280);
INTERCONNECT Split_351_n744_AND2T_122_n161(net281_c1,net281);
INTERCONNECT Split_288_n681_Split_289_n682(net282_c1,net282);
INTERCONNECT Split_264_n657_DFFT_166__FPB_n559(net283_c1,net283);
INTERCONNECT Split_272_n665_OR2T_63_n87(net284_c1,net284);
INTERCONNECT Split_280_n673_AND2T_90_n114(net285_c1,net285);
INTERCONNECT Split_336_n729_Split_337_n730(net286_c1,net286);
INTERCONNECT Split_344_n737_OR2T_105_n129(net287_c1,net287);
INTERCONNECT Split_352_n745_DFFT_234__FPB_n627(net288_c1,net288);
INTERCONNECT Split_360_n753_Split_361_n754(net289_c1,net289);
INTERCONNECT Split_289_n682_AND2T_31_n55(net290_c1,net290);
INTERCONNECT Split_297_n690_AND2T_44_n68(net291_c1,net291);
INTERCONNECT Split_265_n658_DFFT_208__FPB_n601(net292_c1,net292);
INTERCONNECT Split_273_n666_DFFT_153__FPB_n546(net293_c1,net293);
INTERCONNECT Split_281_n674_Split_282_n675(net294_c1,net294);
INTERCONNECT Split_345_n738_DFFT_200__FPB_n593(net295_c1,net295);
INTERCONNECT Split_353_n746_NOTT_119_n158(net296_c1,net296);
INTERCONNECT Split_361_n754_AND2T_17_n41(net297_c1,net297);
INTERCONNECT Split_298_n691_OR2T_46_n70(net298_c1,net298);
INTERCONNECT Split_266_n659_OR2T_82_n106(net299_c1,net299);
INTERCONNECT Split_274_n667_AND2T_79_n103(net300_c1,net300);
INTERCONNECT Split_282_n675_AND2T_25_n49(net301_c1,net301);
INTERCONNECT Split_290_n683_AND2T_79_n103(net302_c1,net302);
INTERCONNECT Split_346_n739_OR2T_105_n129(net303_c1,net303);
INTERCONNECT Split_354_n747_Split_355_n748(net304_c1,net304);
INTERCONNECT Split_362_n755_DFFT_146__FPB_n539(net305_c1,net305);
INTERCONNECT Split_299_n692_Split_300_n693(net306_c1,net306);
INTERCONNECT Split_275_n668_AND2T_88_n112(net307_c1,net307);
INTERCONNECT Split_283_n676_OR2T_76_n100(net308_c1,net308);
INTERCONNECT Split_291_n684_DFFT_221__FPB_n614(net309_c1,net309);
INTERCONNECT Split_355_n748_NOTT_11_n35(net310_c1,net310);
INTERCONNECT Split_363_n756_Split_364_n757(net311_c1,net311);
INTERCONNECT Split_276_n669_DFFT_175__FPB_n568(net312_c1,net312);
INTERCONNECT Split_284_n677_AND2T_26_n50(net313_c1,net313);
INTERCONNECT Split_292_n685_AND2T_30_n54(net314_c1,net314);
INTERCONNECT Split_356_n749_DFFT_151__FPB_n544(net315_c1,net315);
INTERCONNECT Split_364_n757_NOTT_9_n33(net316_c1,net316);
INTERCONNECT Split_300_n693_DFFT_133__FBL_n526(net317_c1,net317);
INTERCONNECT Split_285_n678_Split_286_n679(net318_c1,net318);
INTERCONNECT Split_293_n686_OR2T_37_n61(net319_c1,net319);
INTERCONNECT Split_365_n758_OR2T_83_n107(net320_c1,net320);
INTERCONNECT Split_301_n694_DFFT_138__FBL_n531(net321_c1,net321);
INTERCONNECT Split_286_n679_AND2T_98_n122(net322_c1,net322);
INTERCONNECT Split_294_n687_Split_295_n688(net323_c1,net323);
INTERCONNECT Split_302_n695_OR2T_100_n124(net324_c1,net324);
INTERCONNECT Split_295_n688_OR2T_42_n66(net325_c1,net325);
INTERCONNECT Split_303_n696_AND2T_54_n78(net326_c1,net326);
INTERCONNECT Split_296_n689_AND2T_69_n93(net327_c1,net327);
INTERCONNECT Split_304_n697_AND2T_60_n84(net328_c1,net328);
INTERCONNECT Split_305_n698_DFFT_143__FBL_n536(net329_c1,net329);
INTERCONNECT Split_306_n699_DFFT_134__FBL_n527(net330_c1,net330);
INTERCONNECT DFFT_129__PIPL_n180_DFFT_235__FPB_n628(net331_c1,net331);
INTERCONNECT DFFT_130__PIPL_n181_DFFT_242__FPB_n635(net332_c1,net332);
INTERCONNECT DFFT_131__PIPL_n182_DFFT_249__FPB_n642(net333_c1,net333);
INTERCONNECT DFFT_132__PIPL_n183_DFFT_255__FPB_n648(net334_c1,net334);
INTERCONNECT DFFT_137__FBL_n530_NOTT_120_n159(net335_c1,net335);
INTERCONNECT DFFT_138__FBL_n531_Split_347_n740(net336_c1,net336);
INTERCONNECT DFFT_139__FBL_n532_NOTT_121_n160(net337_c1,net337);
INTERCONNECT DFFT_140__FBL_n533_Split_350_n743(net338_c1,net338);
INTERCONNECT DFFT_141__FBL_n534_Split_352_n745(net339_c1,net339);
INTERCONNECT DFFT_133__FBL_n526_Split_339_n732(net340_c1,net340);
INTERCONNECT DFFT_142__FBL_n535_Split_354_n747(net341_c1,net341);
INTERCONNECT DFFT_134__FBL_n527_Split_340_n733(net342_c1,net342);
INTERCONNECT DFFT_143__FBL_n536_Split_357_n750(net343_c1,net343);
INTERCONNECT DFFT_135__FBL_n528_Split_343_n736(net344_c1,net344);
INTERCONNECT DFFT_144__FBL_n537_Split_360_n753(net345_c1,net345);
INTERCONNECT DFFT_136__FBL_n529_Split_346_n739(net346_c1,net346);
INTERCONNECT DFFT_145__FBL_n538_Split_363_n756(net347_c1,net347);
INTERCONNECT DFFT_207__FPB_n600_OR2T_94_n118(net348_c1,net348);
INTERCONNECT DFFT_208__FPB_n601_DFFT_209__FPB_n602(net349_c1,net349);
INTERCONNECT DFFT_217__FPB_n610_DFFT_218__FPB_n611(net350_c1,net350);
INTERCONNECT DFFT_209__FPB_n602_DFFT_210__FPB_n603(net351_c1,net351);
INTERCONNECT DFFT_127__FPB_n178_Split_333_n726(net352_c1,net352);
INTERCONNECT DFFT_218__FPB_n611_DFFT_219__FPB_n612(net353_c1,net353);
INTERCONNECT DFFT_210__FPB_n603_DFFT_211__FPB_n604(net354_c1,net354);
INTERCONNECT DFFT_128__FPB_n179_Split_336_n729(net355_c1,net355);
INTERCONNECT DFFT_227__FPB_n620_DFFT_228__FPB_n621(net356_c1,net356);
INTERCONNECT DFFT_211__FPB_n604_DFFT_212__FPB_n605(net357_c1,net357);
INTERCONNECT DFFT_219__FPB_n612_AND2T_101_n125(net358_c1,net358);
INTERCONNECT DFFT_147__FPB_n540_AND2T_12_n36(net359_c1,net359);
INTERCONNECT DFFT_228__FPB_n621_DFFT_229__FPB_n622(net360_c1,net360);
INTERCONNECT DFFT_212__FPB_n605_DFFT_213__FPB_n606(net361_c1,net361);
INTERCONNECT DFFT_220__FPB_n613_AND2T_102_n126(net362_c1,net362);
INTERCONNECT DFFT_148__FPB_n541_AND2T_13_n37(net363_c1,net363);
INTERCONNECT DFFT_237__FPB_n630_DFFT_238__FPB_n631(net364_c1,net364);
INTERCONNECT DFFT_229__FPB_n622_DFFT_230__FPB_n623(net365_c1,net365);
INTERCONNECT DFFT_221__FPB_n614_AND2T_103_n127(net366_c1,net366);
INTERCONNECT DFFT_213__FPB_n606_AND2T_95_n119(net367_c1,net367);
INTERCONNECT DFFT_157__FPB_n550_AND2T_34_n58(net368_c1,net368);
INTERCONNECT DFFT_149__FPB_n542_AND2T_14_n38(net369_c1,net369);
INTERCONNECT DFFT_238__FPB_n631_DFFT_239__FPB_n632(net370_c1,net370);
INTERCONNECT DFFT_230__FPB_n623_DFFT_231__FPB_n624(net371_c1,net371);
INTERCONNECT DFFT_214__FPB_n607_DFFT_215__FPB_n608(net372_c1,net372);
INTERCONNECT DFFT_222__FPB_n615_OR2T_106_n130(net373_c1,net373);
INTERCONNECT DFFT_158__FPB_n551_OR2T_37_n61(net374_c1,net374);
INTERCONNECT DFFT_150__FPB_n543_AND2T_16_n40(net375_c1,net375);
INTERCONNECT DFFT_247__FPB_n640_DFFT_248_state_obs1(net376_c1,net376);
INTERCONNECT DFFT_239__FPB_n632_DFFT_240__FPB_n633(net377_c1,net377);
INTERCONNECT DFFT_231__FPB_n624_DFFT_232__FPB_n625(net378_c1,net378);
INTERCONNECT DFFT_167__FPB_n560_DFFT_168__FPB_n561(net379_c1,net379);
INTERCONNECT DFFT_159__FPB_n552_DFFT_160__FPB_n553(net380_c1,net380);
INTERCONNECT DFFT_223__FPB_n616_AND2T_107_n131(net381_c1,net381);
INTERCONNECT DFFT_215__FPB_n608_OR2T_99_n123(net382_c1,net382);
INTERCONNECT DFFT_151__FPB_n544_AND2T_19_n43(net383_c1,net383);
INTERCONNECT DFFT_240__FPB_n633_DFFT_241_state_obs0(net384_c1,net384);
INTERCONNECT DFFT_216__FPB_n609_Split_HOLD_621(net385_c1,net385);
INTERCONNECT DFFT_168__FPB_n561_DFFT_169__FPB_n562(net386_c1,net386);
INTERCONNECT DFFT_160__FPB_n553_DFFT_161__FPB_n554(net387_c1,net387);
INTERCONNECT DFFT_232__FPB_n625_AND2T_114_n138(net388_c1,net388);
INTERCONNECT DFFT_224__FPB_n617_AND2T_109_n133(net389_c1,net389);
INTERCONNECT DFFT_152__FPB_n545_AND2T_20_n44(net390_c1,net390);
INTERCONNECT DFFT_257__FPB_n650_DFFT_258__FPB_n651(net391_c1,net391);
INTERCONNECT DFFT_249__FPB_n642_DFFT_250__FPB_n643(net392_c1,net392);
INTERCONNECT DFFT_169__FPB_n562_DFFT_170__FPB_n563(net393_c1,net393);
INTERCONNECT DFFT_233__FPB_n626_OR2T_116_n140(net394_c1,net394);
INTERCONNECT DFFT_225__FPB_n618_AND2T_110_n134(net395_c1,net395);
INTERCONNECT DFFT_177__FPB_n570_AND2T_59_n83(net396_c1,net396);
INTERCONNECT DFFT_161__FPB_n554_AND2T_38_n62(net397_c1,net397);
INTERCONNECT DFFT_153__FPB_n546_AND2T_21_n45(net398_c1,net398);
INTERCONNECT DFFT_258__FPB_n651_DFFT_259_state_obs3(net399_c1,net399);
INTERCONNECT DFFT_250__FPB_n643_DFFT_251__FPB_n644(net400_c1,net400);
INTERCONNECT DFFT_242__FPB_n635_DFFT_243__FPB_n636(net401_c1,net401);
INTERCONNECT DFFT_170__FPB_n563_DFFT_171__FPB_n564(net402_c1,net402);
INTERCONNECT DFFT_234__FPB_n627_AND2T_125_n164(net403_c1,net403);
INTERCONNECT DFFT_226__FPB_n619_OR2T_112_n136(net404_c1,net404);
INTERCONNECT DFFT_178__FPB_n571_AND2T_60_n84(net405_c1,net405);
INTERCONNECT DFFT_162__FPB_n555_AND2T_39_n63(net406_c1,net406);
INTERCONNECT DFFT_154__FPB_n547_OR2T_23_n47(net407_c1,net407);
INTERCONNECT DFFT_146__FPB_n539_AND2T_10_n34(net408_c1,net408);
INTERCONNECT DFFT_251__FPB_n644_DFFT_252__FPB_n645(net409_c1,net409);
INTERCONNECT DFFT_243__FPB_n636_DFFT_244__FPB_n637(net410_c1,net410);
INTERCONNECT DFFT_235__FPB_n628_DFFT_236__FPB_n629(net411_c1,net411);
INTERCONNECT DFFT_187__FPB_n580_AND2T_69_n93(net412_c1,net412);
INTERCONNECT DFFT_179__FPB_n572_OR2T_63_n87(net413_c1,net413);
INTERCONNECT DFFT_171__FPB_n564_AND2T_50_n74(net414_c1,net414);
INTERCONNECT DFFT_163__FPB_n556_AND2T_41_n65(net415_c1,net415);
INTERCONNECT DFFT_155__FPB_n548_AND2T_26_n50(net416_c1,net416);
INTERCONNECT DFFT_252__FPB_n645_DFFT_253__FPB_n646(net417_c1,net417);
INTERCONNECT DFFT_244__FPB_n637_DFFT_245__FPB_n638(net418_c1,net418);
INTERCONNECT DFFT_236__FPB_n629_DFFT_237__FPB_n630(net419_c1,net419);
INTERCONNECT DFFT_188__FPB_n581_DFFT_189__FPB_n582(net420_c1,net420);
INTERCONNECT DFFT_180__FPB_n573_AND2T_64_n88(net421_c1,net421);
INTERCONNECT DFFT_172__FPB_n565_AND2T_51_n75(net422_c1,net422);
INTERCONNECT DFFT_164__FPB_n557_AND2T_43_n67(net423_c1,net423);
INTERCONNECT DFFT_156__FPB_n549_OR2T_32_n56(net424_c1,net424);
INTERCONNECT DFFT_253__FPB_n646_DFFT_254_state_obs2(net425_c1,net425);
INTERCONNECT DFFT_245__FPB_n638_DFFT_246__FPB_n639(net426_c1,net426);
INTERCONNECT DFFT_197__FPB_n590_DFFT_198__FPB_n591(net427_c1,net427);
INTERCONNECT DFFT_189__FPB_n582_DFFT_190__FPB_n583(net428_c1,net428);
INTERCONNECT DFFT_181__FPB_n574_DFFT_182__FPB_n575(net429_c1,net429);
INTERCONNECT DFFT_173__FPB_n566_DFFT_174__FPB_n567(net430_c1,net430);
INTERCONNECT DFFT_165__FPB_n558_OR2T_46_n70(net431_c1,net431);
INTERCONNECT DFFT_246__FPB_n639_DFFT_247__FPB_n640(net432_c1,net432);
INTERCONNECT DFFT_198__FPB_n591_DFFT_199__FPB_n592(net433_c1,net433);
INTERCONNECT DFFT_190__FPB_n583_DFFT_191__FPB_n584(net434_c1,net434);
INTERCONNECT DFFT_182__FPB_n575_DFFT_183__FPB_n576(net435_c1,net435);
INTERCONNECT DFFT_166__FPB_n559_DFFT_167__FPB_n560(net436_c1,net436);
INTERCONNECT DFFT_174__FPB_n567_AND2T_54_n78(net437_c1,net437);
INTERCONNECT DFFT_255__FPB_n648_DFFT_256__FPB_n649(net438_c1,net438);
INTERCONNECT DFFT_191__FPB_n584_DFFT_192__FPB_n585(net439_c1,net439);
INTERCONNECT DFFT_199__FPB_n592_AND2T_78_n102(net440_c1,net440);
INTERCONNECT DFFT_183__FPB_n576_AND2T_66_n90(net441_c1,net441);
INTERCONNECT DFFT_175__FPB_n568_AND2T_56_n80(net442_c1,net442);
INTERCONNECT DFFT_256__FPB_n649_DFFT_257__FPB_n650(net443_c1,net443);
INTERCONNECT DFFT_200__FPB_n593_DFFT_201__FPB_n594(net444_c1,net444);
INTERCONNECT DFFT_192__FPB_n585_DFFT_193__FPB_n586(net445_c1,net445);
INTERCONNECT DFFT_184__FPB_n577_DFFT_185__FPB_n578(net446_c1,net446);
INTERCONNECT DFFT_176__FPB_n569_AND2T_58_n82(net447_c1,net447);
INTERCONNECT DFFT_201__FPB_n594_AND2T_81_n105(net448_c1,net448);
INTERCONNECT DFFT_193__FPB_n586_AND2T_74_n98(net449_c1,net449);
INTERCONNECT DFFT_185__FPB_n578_AND2T_67_n91(net450_c1,net450);
INTERCONNECT DFFT_186__FPB_n579_DFFT_187__FPB_n580(net451_c1,net451);
INTERCONNECT DFFT_202__FPB_n595_AND2T_84_n108(net452_c1,net452);
INTERCONNECT DFFT_194__FPB_n587_OR2T_75_n99(net453_c1,net453);
INTERCONNECT DFFT_203__FPB_n596_AND2T_85_n109(net454_c1,net454);
INTERCONNECT DFFT_195__FPB_n588_OR2T_76_n100(net455_c1,net455);
INTERCONNECT DFFT_204__FPB_n597_AND2T_86_n110(net456_c1,net456);
INTERCONNECT DFFT_196__FPB_n589_AND2T_77_n101(net457_c1,net457);
INTERCONNECT DFFT_205__FPB_n598_AND2T_91_n115(net458_c1,net458);
INTERCONNECT DFFT_206__FPB_n599_OR2T_93_n117(net459_c1,net459);
INTERCONNECT DFFT_241_state_obs0_state_obs0_Pad(net460_c1,state_obs0_Pad);
INTERCONNECT DFFT_248_state_obs1_state_obs1_Pad(net461_c1,state_obs1_Pad);
INTERCONNECT DFFT_254_state_obs2_state_obs2_Pad(net462_c1,state_obs2_Pad);
INTERCONNECT DFFT_259_state_obs3_state_obs3_Pad(net463_c1,state_obs3_Pad);
INTERCONNECT DFFT_117_state0_buf_DFFT_129__PIPL_n180(net464_c1,net464);
INTERCONNECT DFFT_118_state1_buf_DFFT_130__PIPL_n181(net465_c1,net465);
INTERCONNECT SplitCLK_0_507_SplitCLK_0_377(net466_c1,net466);
INTERCONNECT SplitCLK_0_507_SplitCLK_2_502(net467_c1,net467);
INTERCONNECT SplitCLK_2_506_DFFT_169__FPB_n562(net468_c1,net468);
INTERCONNECT SplitCLK_2_505_DFFT_182__FPB_n575(net469_c1,net469);
INTERCONNECT SplitCLK_2_504_DFFT_229__FPB_n622(net470_c1,net470);
INTERCONNECT SplitCLK_2_503_DFFT_225__FPB_n618(net471_c1,net471);
INTERCONNECT SplitCLK_2_502_SplitCLK_6_439(net472_c1,net472);
INTERCONNECT SplitCLK_2_502_SplitCLK_4_501(net473_c1,net473);
INTERCONNECT SplitCLK_4_501_SplitCLK_4_470(net474_c1,net474);
INTERCONNECT SplitCLK_4_501_SplitCLK_2_500(net475_c1,net475);
INTERCONNECT SplitCLK_2_500_SplitCLK_6_485(net476_c1,net476);
INTERCONNECT SplitCLK_2_500_SplitCLK_4_499(net477_c1,net477);
INTERCONNECT SplitCLK_4_499_SplitCLK_4_492(net478_c1,net478);
INTERCONNECT SplitCLK_4_499_SplitCLK_2_498(net479_c1,net479);
INTERCONNECT SplitCLK_2_498_SplitCLK_2_495(net480_c1,net480);
INTERCONNECT SplitCLK_2_498_SplitCLK_2_497(net481_c1,net481);
INTERCONNECT SplitCLK_2_497_SplitCLK_2_506(net482_c1,net482);
INTERCONNECT SplitCLK_2_497_SplitCLK_4_496(net483_c1,net483);
INTERCONNECT SplitCLK_4_496_DFFT_170__FPB_n563(net484_c1,net484);
INTERCONNECT SplitCLK_4_496_DFFT_168__FPB_n561(net485_c1,net485);
INTERCONNECT SplitCLK_2_495_SplitCLK_4_493(net486_c1,net486);
INTERCONNECT SplitCLK_2_495_SplitCLK_4_494(net487_c1,net487);
INTERCONNECT SplitCLK_4_494_DFFT_142__FBL_n535(net488_c1,net488);
INTERCONNECT SplitCLK_4_494_DFFT_158__FPB_n551(net489_c1,net489);
INTERCONNECT SplitCLK_4_493_OR2T_37_n61(net490_c1,net490);
INTERCONNECT SplitCLK_4_493_DFFT_171__FPB_n564(net491_c1,net491);
INTERCONNECT SplitCLK_4_492_SplitCLK_4_488(net492_c1,net492);
INTERCONNECT SplitCLK_4_492_SplitCLK_4_491(net493_c1,net493);
INTERCONNECT SplitCLK_4_491_SplitCLK_4_489(net494_c1,net494);
INTERCONNECT SplitCLK_4_491_SplitCLK_2_490(net495_c1,net495);
INTERCONNECT SplitCLK_2_490_AND2T_50_n74(net496_c1,net496);
INTERCONNECT SplitCLK_2_490_DFFT_167__FPB_n560(net497_c1,net497);
INTERCONNECT SplitCLK_4_489_DFFT_166__FPB_n559(net498_c1,net498);
INTERCONNECT SplitCLK_4_489_DFFT_188__FPB_n581(net499_c1,net499);
INTERCONNECT SplitCLK_4_488_SplitCLK_4_486(net500_c1,net500);
INTERCONNECT SplitCLK_4_488_SplitCLK_4_487(net501_c1,net501);
INTERCONNECT SplitCLK_4_487_AND2T_36_n60(net502_c1,net502);
INTERCONNECT SplitCLK_4_487_DFFT_137__FBL_n530(net503_c1,net503);
INTERCONNECT SplitCLK_4_486_DFFT_154__FPB_n547(net504_c1,net504);
INTERCONNECT SplitCLK_4_486_NOTT_120_n159(net505_c1,net505);
INTERCONNECT SplitCLK_6_485_SplitCLK_0_477(net506_c1,net506);
INTERCONNECT SplitCLK_6_485_SplitCLK_2_484(net507_c1,net507);
INTERCONNECT SplitCLK_2_484_SplitCLK_6_480(net508_c1,net508);
INTERCONNECT SplitCLK_2_484_SplitCLK_4_483(net509_c1,net509);
INTERCONNECT SplitCLK_4_483_SplitCLK_4_481(net510_c1,net510);
INTERCONNECT SplitCLK_4_483_SplitCLK_4_482(net511_c1,net511);
INTERCONNECT SplitCLK_4_482_AND2T_64_n88(net512_c1,net512);
INTERCONNECT SplitCLK_4_482_DFFT_180__FPB_n573(net513_c1,net513);
INTERCONNECT SplitCLK_4_481_OR2T_65_n89(net514_c1,net514);
INTERCONNECT SplitCLK_4_481_DFFT_152__FPB_n545(net515_c1,net515);
INTERCONNECT SplitCLK_6_480_SplitCLK_4_478(net516_c1,net516);
INTERCONNECT SplitCLK_6_480_SplitCLK_4_479(net517_c1,net517);
INTERCONNECT SplitCLK_4_479_OR2T_63_n87(net518_c1,net518);
INTERCONNECT SplitCLK_4_479_DFFT_179__FPB_n572(net519_c1,net519);
INTERCONNECT SplitCLK_4_478_AND2T_66_n90(net520_c1,net520);
INTERCONNECT SplitCLK_4_478_DFFT_138__FBL_n531(net521_c1,net521);
INTERCONNECT SplitCLK_0_477_SplitCLK_6_473(net522_c1,net522);
INTERCONNECT SplitCLK_0_477_SplitCLK_0_476(net523_c1,net523);
INTERCONNECT SplitCLK_0_476_SplitCLK_4_474(net524_c1,net524);
INTERCONNECT SplitCLK_0_476_SplitCLK_0_475(net525_c1,net525);
INTERCONNECT SplitCLK_0_475_DFFT_139__FBL_n532(net526_c1,net526);
INTERCONNECT SplitCLK_0_475_NOTT_121_n160(net527_c1,net527);
INTERCONNECT SplitCLK_4_474_DFFT_143__FBL_n536(net528_c1,net528);
INTERCONNECT SplitCLK_4_474_DFFT_151__FPB_n544(net529_c1,net529);
INTERCONNECT SplitCLK_6_473_SplitCLK_4_471(net530_c1,net530);
INTERCONNECT SplitCLK_6_473_SplitCLK_4_472(net531_c1,net531);
INTERCONNECT SplitCLK_4_472_OR2T_72_n96(net532_c1,net532);
INTERCONNECT SplitCLK_4_472_DFFT_183__FPB_n576(net533_c1,net533);
INTERCONNECT SplitCLK_4_471_OR2T_73_n97(net534_c1,net534);
INTERCONNECT SplitCLK_4_471_DFFT_134__FBL_n527(net535_c1,net535);
INTERCONNECT SplitCLK_4_470_SplitCLK_2_454(net536_c1,net536);
INTERCONNECT SplitCLK_4_470_SplitCLK_4_469(net537_c1,net537);
INTERCONNECT SplitCLK_4_469_SplitCLK_0_461(net538_c1,net538);
INTERCONNECT SplitCLK_4_469_SplitCLK_6_468(net539_c1,net539);
INTERCONNECT SplitCLK_6_468_SplitCLK_4_464(net540_c1,net540);
INTERCONNECT SplitCLK_6_468_SplitCLK_4_467(net541_c1,net541);
INTERCONNECT SplitCLK_4_467_SplitCLK_4_465(net542_c1,net542);
INTERCONNECT SplitCLK_4_467_SplitCLK_4_466(net543_c1,net543);
INTERCONNECT SplitCLK_4_466_DFFT_190__FPB_n583(net544_c1,net544);
INTERCONNECT SplitCLK_4_466_DFFT_189__FPB_n582(net545_c1,net545);
INTERCONNECT SplitCLK_4_465_DFFT_191__FPB_n584(net546_c1,net546);
INTERCONNECT SplitCLK_4_465_DFFT_193__FPB_n586(net547_c1,net547);
INTERCONNECT SplitCLK_4_464_SplitCLK_4_462(net548_c1,net548);
INTERCONNECT SplitCLK_4_464_SplitCLK_0_463(net549_c1,net549);
INTERCONNECT SplitCLK_0_463_AND2T_45_n69(net550_c1,net550);
INTERCONNECT SplitCLK_0_463_OR2T_23_n47(net551_c1,net551);
INTERCONNECT SplitCLK_4_462_NOTT_123_n162(net552_c1,net552);
INTERCONNECT SplitCLK_4_462_DFFT_176__FPB_n569(net553_c1,net553);
INTERCONNECT SplitCLK_0_461_SplitCLK_6_457(net554_c1,net554);
INTERCONNECT SplitCLK_0_461_SplitCLK_4_460(net555_c1,net555);
INTERCONNECT SplitCLK_4_460_SplitCLK_4_458(net556_c1,net556);
INTERCONNECT SplitCLK_4_460_SplitCLK_4_459(net557_c1,net557);
INTERCONNECT SplitCLK_4_459_DFFT_155__FPB_n548(net558_c1,net558);
INTERCONNECT SplitCLK_4_459_DFFT_192__FPB_n585(net559_c1,net559);
INTERCONNECT SplitCLK_4_458_DFFT_230__FPB_n623(net560_c1,net560);
INTERCONNECT SplitCLK_4_458_DFFT_231__FPB_n624(net561_c1,net561);
INTERCONNECT SplitCLK_6_457_SplitCLK_4_455(net562_c1,net562);
INTERCONNECT SplitCLK_6_457_SplitCLK_4_456(net563_c1,net563);
INTERCONNECT SplitCLK_4_456_AND2T_30_n54(net564_c1,net564);
INTERCONNECT SplitCLK_4_456_OR2T_46_n70(net565_c1,net565);
INTERCONNECT SplitCLK_4_455_AND2T_26_n50(net566_c1,net566);
INTERCONNECT SplitCLK_4_455_AND2T_19_n43(net567_c1,net567);
INTERCONNECT SplitCLK_2_454_SplitCLK_4_446(net568_c1,net568);
INTERCONNECT SplitCLK_2_454_SplitCLK_6_453(net569_c1,net569);
INTERCONNECT SplitCLK_6_453_SplitCLK_6_449(net570_c1,net570);
INTERCONNECT SplitCLK_6_453_SplitCLK_6_452(net571_c1,net571);
INTERCONNECT SplitCLK_6_452_SplitCLK_4_450(net572_c1,net572);
INTERCONNECT SplitCLK_6_452_SplitCLK_4_451(net573_c1,net573);
INTERCONNECT SplitCLK_4_451_AND2T_43_n67(net574_c1,net574);
INTERCONNECT SplitCLK_4_451_AND2T_74_n98(net575_c1,net575);
INTERCONNECT SplitCLK_4_450_AND2T_35_n59(net576_c1,net576);
INTERCONNECT SplitCLK_4_450_NOTT_15_n39(net577_c1,net577);
INTERCONNECT SplitCLK_6_449_SplitCLK_4_447(net578_c1,net578);
INTERCONNECT SplitCLK_6_449_SplitCLK_4_448(net579_c1,net579);
INTERCONNECT SplitCLK_4_448_OR2T_71_n95(net580_c1,net580);
INTERCONNECT SplitCLK_4_448_DFFT_164__FPB_n557(net581_c1,net581);
INTERCONNECT SplitCLK_4_447_AND2T_68_n92(net582_c1,net582);
INTERCONNECT SplitCLK_4_447_OR2T_70_n94(net583_c1,net583);
INTERCONNECT SplitCLK_4_446_SplitCLK_6_442(net584_c1,net584);
INTERCONNECT SplitCLK_4_446_SplitCLK_4_445(net585_c1,net585);
INTERCONNECT SplitCLK_4_445_SplitCLK_4_443(net586_c1,net586);
INTERCONNECT SplitCLK_4_445_SplitCLK_4_444(net587_c1,net587);
INTERCONNECT SplitCLK_4_444_AND2T_44_n68(net588_c1,net588);
INTERCONNECT SplitCLK_4_444_DFFT_165__FPB_n558(net589_c1,net589);
INTERCONNECT SplitCLK_4_443_AND2T_58_n82(net590_c1,net590);
INTERCONNECT SplitCLK_4_443_OR2T_89_n113(net591_c1,net591);
INTERCONNECT SplitCLK_6_442_SplitCLK_4_440(net592_c1,net592);
INTERCONNECT SplitCLK_6_442_SplitCLK_4_441(net593_c1,net593);
INTERCONNECT SplitCLK_4_441_OR2T_57_n81(net594_c1,net594);
INTERCONNECT SplitCLK_4_441_AND2T_90_n114(net595_c1,net595);
INTERCONNECT SplitCLK_4_440_OR2T_61_n85(net596_c1,net596);
INTERCONNECT SplitCLK_4_440_OR2T_62_n86(net597_c1,net597);
INTERCONNECT SplitCLK_6_439_SplitCLK_0_408(net598_c1,net598);
INTERCONNECT SplitCLK_6_439_SplitCLK_6_438(net599_c1,net599);
INTERCONNECT SplitCLK_6_438_SplitCLK_6_423(net600_c1,net600);
INTERCONNECT SplitCLK_6_438_SplitCLK_4_437(net601_c1,net601);
INTERCONNECT SplitCLK_4_437_SplitCLK_0_430(net602_c1,net602);
INTERCONNECT SplitCLK_4_437_SplitCLK_4_436(net603_c1,net603);
INTERCONNECT SplitCLK_4_436_SplitCLK_0_433(net604_c1,net604);
INTERCONNECT SplitCLK_4_436_SplitCLK_2_435(net605_c1,net605);
INTERCONNECT SplitCLK_2_435_SplitCLK_2_505(net606_c1,net606);
INTERCONNECT SplitCLK_2_435_SplitCLK_4_434(net607_c1,net607);
INTERCONNECT SplitCLK_4_434_AND2T_51_n75(net608_c1,net608);
INTERCONNECT SplitCLK_4_434_DFFT_172__FPB_n565(net609_c1,net609);
INTERCONNECT SplitCLK_0_433_SplitCLK_4_431(net610_c1,net610);
INTERCONNECT SplitCLK_0_433_SplitCLK_0_432(net611_c1,net611);
INTERCONNECT SplitCLK_0_432_AND2T_84_n108(net612_c1,net612);
INTERCONNECT SplitCLK_0_432_DFFT_173__FPB_n566(net613_c1,net613);
INTERCONNECT SplitCLK_4_431_AND2T_85_n109(net614_c1,net614);
INTERCONNECT SplitCLK_4_431_DFFT_174__FPB_n567(net615_c1,net615);
INTERCONNECT SplitCLK_0_430_SplitCLK_6_426(net616_c1,net616);
INTERCONNECT SplitCLK_0_430_SplitCLK_4_429(net617_c1,net617);
INTERCONNECT SplitCLK_4_429_SplitCLK_4_427(net618_c1,net618);
INTERCONNECT SplitCLK_4_429_SplitCLK_4_428(net619_c1,net619);
INTERCONNECT SplitCLK_4_428_AND2T_28_n52(net620_c1,net620);
INTERCONNECT SplitCLK_4_428_DFFT_202__FPB_n595(net621_c1,net621);
INTERCONNECT SplitCLK_4_427_AND2T_122_n161(net622_c1,net622);
INTERCONNECT SplitCLK_4_427_NOTT_126_n177(net623_c1,net623);
INTERCONNECT SplitCLK_6_426_SplitCLK_4_424(net624_c1,net624);
INTERCONNECT SplitCLK_6_426_SplitCLK_4_425(net625_c1,net625);
INTERCONNECT SplitCLK_4_425_DFFT_203__FPB_n596(net626_c1,net626);
INTERCONNECT SplitCLK_4_425_OR2T_83_n107(net627_c1,net627);
INTERCONNECT SplitCLK_4_424_AND2T_86_n110(net628_c1,net628);
INTERCONNECT SplitCLK_4_424_DFFT_204__FPB_n597(net629_c1,net629);
INTERCONNECT SplitCLK_6_423_SplitCLK_6_415(net630_c1,net630);
INTERCONNECT SplitCLK_6_423_SplitCLK_6_422(net631_c1,net631);
INTERCONNECT SplitCLK_6_422_SplitCLK_6_418(net632_c1,net632);
INTERCONNECT SplitCLK_6_422_SplitCLK_6_421(net633_c1,net633);
INTERCONNECT SplitCLK_6_421_SplitCLK_4_419(net634_c1,net634);
INTERCONNECT SplitCLK_6_421_SplitCLK_4_420(net635_c1,net635);
INTERCONNECT SplitCLK_4_420_DFFT_117_state0_buf(net636_c1,net636);
INTERCONNECT SplitCLK_4_420_DFFT_181__FPB_n574(net637_c1,net637);
INTERCONNECT SplitCLK_4_419_DFFT_129__PIPL_n180(net638_c1,net638);
INTERCONNECT SplitCLK_4_419_DFFT_128__FPB_n179(net639_c1,net639);
INTERCONNECT SplitCLK_6_418_SplitCLK_4_416(net640_c1,net640);
INTERCONNECT SplitCLK_6_418_SplitCLK_0_417(net641_c1,net641);
INTERCONNECT SplitCLK_0_417_DFFT_241_state_obs0(net642_c1,net642);
INTERCONNECT SplitCLK_0_417_DFFT_240__FPB_n633(net643_c1,net643);
INTERCONNECT SplitCLK_4_416_DFFT_235__FPB_n628(net644_c1,net644);
INTERCONNECT SplitCLK_4_416_DFFT_239__FPB_n632(net645_c1,net645);
INTERCONNECT SplitCLK_6_415_SplitCLK_6_411(net646_c1,net646);
INTERCONNECT SplitCLK_6_415_SplitCLK_2_414(net647_c1,net647);
INTERCONNECT SplitCLK_2_414_SplitCLK_4_412(net648_c1,net648);
INTERCONNECT SplitCLK_2_414_SplitCLK_4_413(net649_c1,net649);
INTERCONNECT SplitCLK_4_413_DFFT_222__FPB_n615(net650_c1,net650);
INTERCONNECT SplitCLK_4_413_OR2T_82_n106(net651_c1,net651);
INTERCONNECT SplitCLK_4_412_DFFT_133__FBL_n526(net652_c1,net652);
INTERCONNECT SplitCLK_4_412_DFFT_157__FPB_n550(net653_c1,net653);
INTERCONNECT SplitCLK_6_411_SplitCLK_4_409(net654_c1,net654);
INTERCONNECT SplitCLK_6_411_SplitCLK_4_410(net655_c1,net655);
INTERCONNECT SplitCLK_4_410_DFFT_236__FPB_n629(net656_c1,net656);
INTERCONNECT SplitCLK_4_410_DFFT_237__FPB_n630(net657_c1,net657);
INTERCONNECT SplitCLK_4_409_OR2T_87_n111(net658_c1,net658);
INTERCONNECT SplitCLK_4_409_DFFT_238__FPB_n631(net659_c1,net659);
INTERCONNECT SplitCLK_0_408_SplitCLK_6_392(net660_c1,net660);
INTERCONNECT SplitCLK_0_408_SplitCLK_4_407(net661_c1,net661);
INTERCONNECT SplitCLK_4_407_SplitCLK_0_399(net662_c1,net662);
INTERCONNECT SplitCLK_4_407_SplitCLK_6_406(net663_c1,net663);
INTERCONNECT SplitCLK_6_406_SplitCLK_4_402(net664_c1,net664);
INTERCONNECT SplitCLK_6_406_SplitCLK_4_405(net665_c1,net665);
INTERCONNECT SplitCLK_4_405_SplitCLK_4_403(net666_c1,net666);
INTERCONNECT SplitCLK_4_405_SplitCLK_4_404(net667_c1,net667);
INTERCONNECT SplitCLK_4_404_AND2T_29_n53(net668_c1,net668);
INTERCONNECT SplitCLK_4_404_NOTT_124_n163(net669_c1,net669);
INTERCONNECT SplitCLK_4_403_AND2T_52_n76(net670_c1,net670);
INTERCONNECT SplitCLK_4_403_DFFT_195__FPB_n588(net671_c1,net671);
INTERCONNECT SplitCLK_4_402_SplitCLK_4_400(net672_c1,net672);
INTERCONNECT SplitCLK_4_402_SplitCLK_4_401(net673_c1,net673);
INTERCONNECT SplitCLK_4_401_AND2T_125_n164(net674_c1,net674);
INTERCONNECT SplitCLK_4_401_DFFT_141__FBL_n534(net675_c1,net675);
INTERCONNECT SplitCLK_4_400_OR2T_92_n116(net676_c1,net676);
INTERCONNECT SplitCLK_4_400_DFFT_234__FPB_n627(net677_c1,net677);
INTERCONNECT SplitCLK_0_399_SplitCLK_2_395(net678_c1,net678);
INTERCONNECT SplitCLK_0_399_SplitCLK_4_398(net679_c1,net679);
INTERCONNECT SplitCLK_4_398_SplitCLK_4_396(net680_c1,net680);
INTERCONNECT SplitCLK_4_398_SplitCLK_4_397(net681_c1,net681);
INTERCONNECT SplitCLK_4_397_AND2T_54_n78(net682_c1,net682);
INTERCONNECT SplitCLK_4_397_NOTT_119_n158(net683_c1,net683);
INTERCONNECT SplitCLK_4_396_AND2T_10_n34(net684_c1,net684);
INTERCONNECT SplitCLK_4_396_DFFT_224__FPB_n617(net685_c1,net685);
INTERCONNECT SplitCLK_2_395_SplitCLK_4_393(net686_c1,net686);
INTERCONNECT SplitCLK_2_395_SplitCLK_4_394(net687_c1,net687);
INTERCONNECT SplitCLK_4_394_AND2T_91_n115(net688_c1,net688);
INTERCONNECT SplitCLK_4_394_OR2T_99_n123(net689_c1,net689);
INTERCONNECT SplitCLK_4_393_AND2T_114_n138(net690_c1,net690);
INTERCONNECT SplitCLK_4_393_AND2T_53_n77(net691_c1,net691);
INTERCONNECT SplitCLK_6_392_SplitCLK_0_384(net692_c1,net692);
INTERCONNECT SplitCLK_6_392_SplitCLK_2_391(net693_c1,net693);
INTERCONNECT SplitCLK_2_391_SplitCLK_6_387(net694_c1,net694);
INTERCONNECT SplitCLK_2_391_SplitCLK_2_390(net695_c1,net695);
INTERCONNECT SplitCLK_2_390_SplitCLK_4_388(net696_c1,net696);
INTERCONNECT SplitCLK_2_390_SplitCLK_4_389(net697_c1,net697);
INTERCONNECT SplitCLK_4_389_AND2T_34_n58(net698_c1,net698);
INTERCONNECT SplitCLK_4_389_DFFT_118_state1_buf(net699_c1,net699);
INTERCONNECT SplitCLK_4_388_DFFT_221__FPB_n614(net700_c1,net700);
INTERCONNECT SplitCLK_4_388_DFFT_145__FBL_n538(net701_c1,net701);
INTERCONNECT SplitCLK_6_387_SplitCLK_4_385(net702_c1,net702);
INTERCONNECT SplitCLK_6_387_SplitCLK_4_386(net703_c1,net703);
INTERCONNECT SplitCLK_4_386_DFFT_248_state_obs1(net704_c1,net704);
INTERCONNECT SplitCLK_4_386_DFFT_247__FPB_n640(net705_c1,net705);
INTERCONNECT SplitCLK_4_385_DFFT_130__PIPL_n181(net706_c1,net706);
INTERCONNECT SplitCLK_4_385_DFFT_246__FPB_n639(net707_c1,net707);
INTERCONNECT SplitCLK_0_384_SplitCLK_6_380(net708_c1,net708);
INTERCONNECT SplitCLK_0_384_SplitCLK_4_383(net709_c1,net709);
INTERCONNECT SplitCLK_4_383_SplitCLK_4_381(net710_c1,net710);
INTERCONNECT SplitCLK_4_383_SplitCLK_4_382(net711_c1,net711);
INTERCONNECT SplitCLK_4_382_DFFT_136__FBL_n529(net712_c1,net712);
INTERCONNECT SplitCLK_4_382_DFFT_242__FPB_n635(net713_c1,net713);
INTERCONNECT SplitCLK_4_381_NOTT_9_n33(net714_c1,net714);
INTERCONNECT SplitCLK_4_381_DFFT_205__FPB_n598(net715_c1,net715);
INTERCONNECT SplitCLK_6_380_SplitCLK_4_378(net716_c1,net716);
INTERCONNECT SplitCLK_6_380_SplitCLK_4_379(net717_c1,net717);
INTERCONNECT SplitCLK_4_379_DFFT_244__FPB_n637(net718_c1,net718);
INTERCONNECT SplitCLK_4_379_DFFT_245__FPB_n638(net719_c1,net719);
INTERCONNECT SplitCLK_4_378_AND2T_88_n112(net720_c1,net720);
INTERCONNECT SplitCLK_4_378_DFFT_243__FPB_n636(net721_c1,net721);
INTERCONNECT SplitCLK_0_377_SplitCLK_6_314(net722_c1,net722);
INTERCONNECT SplitCLK_0_377_SplitCLK_4_376(net723_c1,net723);
INTERCONNECT SplitCLK_4_376_SplitCLK_0_345(net724_c1,net724);
INTERCONNECT SplitCLK_4_376_SplitCLK_4_375(net725_c1,net725);
INTERCONNECT SplitCLK_4_375_SplitCLK_6_360(net726_c1,net726);
INTERCONNECT SplitCLK_4_375_SplitCLK_4_374(net727_c1,net727);
INTERCONNECT SplitCLK_4_374_SplitCLK_4_367(net728_c1,net728);
INTERCONNECT SplitCLK_4_374_SplitCLK_6_373(net729_c1,net729);
INTERCONNECT SplitCLK_6_373_SplitCLK_4_370(net730_c1,net730);
INTERCONNECT SplitCLK_6_373_SplitCLK_4_372(net731_c1,net731);
INTERCONNECT SplitCLK_4_372_SplitCLK_2_504(net732_c1,net732);
INTERCONNECT SplitCLK_4_372_SplitCLK_4_371(net733_c1,net733);
INTERCONNECT SplitCLK_4_371_DFFT_227__FPB_n620(net734_c1,net734);
INTERCONNECT SplitCLK_4_371_DFFT_228__FPB_n621(net735_c1,net735);
INTERCONNECT SplitCLK_4_370_SplitCLK_4_368(net736_c1,net736);
INTERCONNECT SplitCLK_4_370_SplitCLK_4_369(net737_c1,net737);
INTERCONNECT SplitCLK_4_369_DFFT_127__FPB_n178(net738_c1,net738);
INTERCONNECT SplitCLK_4_369_DFFT_232__FPB_n625(net739_c1,net739);
INTERCONNECT SplitCLK_4_368_DFFT_156__FPB_n549(net740_c1,net740);
INTERCONNECT SplitCLK_4_368_DFFT_159__FPB_n552(net741_c1,net741);
INTERCONNECT SplitCLK_4_367_SplitCLK_0_363(net742_c1,net742);
INTERCONNECT SplitCLK_4_367_SplitCLK_4_366(net743_c1,net743);
INTERCONNECT SplitCLK_4_366_SplitCLK_4_364(net744_c1,net744);
INTERCONNECT SplitCLK_4_366_SplitCLK_4_365(net745_c1,net745);
INTERCONNECT SplitCLK_4_365_OR2T_33_n57(net746_c1,net746);
INTERCONNECT SplitCLK_4_365_OR2T_49_n73(net747_c1,net747);
INTERCONNECT SplitCLK_4_364_NOTT_8_n32(net748_c1,net748);
INTERCONNECT SplitCLK_4_364_DFFT_208__FPB_n601(net749_c1,net749);
INTERCONNECT SplitCLK_0_363_SplitCLK_4_361(net750_c1,net750);
INTERCONNECT SplitCLK_0_363_SplitCLK_0_362(net751_c1,net751);
INTERCONNECT SplitCLK_0_362_AND2T_31_n55(net752_c1,net752);
INTERCONNECT SplitCLK_0_362_DFFT_149__FPB_n542(net753_c1,net753);
INTERCONNECT SplitCLK_4_361_OR2T_22_n46(net754_c1,net754);
INTERCONNECT SplitCLK_4_361_OR2T_48_n72(net755_c1,net755);
INTERCONNECT SplitCLK_6_360_SplitCLK_6_352(net756_c1,net756);
INTERCONNECT SplitCLK_6_360_SplitCLK_6_359(net757_c1,net757);
INTERCONNECT SplitCLK_6_359_SplitCLK_6_355(net758_c1,net758);
INTERCONNECT SplitCLK_6_359_SplitCLK_2_358(net759_c1,net759);
INTERCONNECT SplitCLK_2_358_SplitCLK_4_356(net760_c1,net760);
INTERCONNECT SplitCLK_2_358_SplitCLK_4_357(net761_c1,net761);
INTERCONNECT SplitCLK_4_357_AND2T_20_n44(net762_c1,net762);
INTERCONNECT SplitCLK_4_357_AND2T_67_n91(net763_c1,net763);
INTERCONNECT SplitCLK_4_356_AND2T_25_n49(net764_c1,net764);
INTERCONNECT SplitCLK_4_356_OR2T_32_n56(net765_c1,net765);
INTERCONNECT SplitCLK_6_355_SplitCLK_4_353(net766_c1,net766);
INTERCONNECT SplitCLK_6_355_SplitCLK_4_354(net767_c1,net767);
INTERCONNECT SplitCLK_4_354_AND2T_109_n133(net768_c1,net768);
INTERCONNECT SplitCLK_4_354_AND2T_60_n84(net769_c1,net769);
INTERCONNECT SplitCLK_4_353_AND2T_59_n83(net770_c1,net770);
INTERCONNECT SplitCLK_4_353_AND2T_69_n93(net771_c1,net771);
INTERCONNECT SplitCLK_6_352_SplitCLK_2_348(net772_c1,net772);
INTERCONNECT SplitCLK_6_352_SplitCLK_4_351(net773_c1,net773);
INTERCONNECT SplitCLK_4_351_SplitCLK_4_349(net774_c1,net774);
INTERCONNECT SplitCLK_4_351_SplitCLK_4_350(net775_c1,net775);
INTERCONNECT SplitCLK_4_350_AND2T_24_n48(net776_c1,net776);
INTERCONNECT SplitCLK_4_350_AND2T_39_n63(net777_c1,net777);
INTERCONNECT SplitCLK_4_349_AND2T_21_n45(net778_c1,net778);
INTERCONNECT SplitCLK_4_349_DFFT_153__FPB_n546(net779_c1,net779);
INTERCONNECT SplitCLK_2_348_SplitCLK_4_346(net780_c1,net780);
INTERCONNECT SplitCLK_2_348_SplitCLK_4_347(net781_c1,net781);
INTERCONNECT SplitCLK_4_347_DFFT_177__FPB_n570(net782_c1,net782);
INTERCONNECT SplitCLK_4_347_DFFT_178__FPB_n571(net783_c1,net783);
INTERCONNECT SplitCLK_4_346_AND2T_40_n64(net784_c1,net784);
INTERCONNECT SplitCLK_4_346_DFFT_187__FPB_n580(net785_c1,net785);
INTERCONNECT SplitCLK_0_345_SplitCLK_6_329(net786_c1,net786);
INTERCONNECT SplitCLK_0_345_SplitCLK_4_344(net787_c1,net787);
INTERCONNECT SplitCLK_4_344_SplitCLK_4_336(net788_c1,net788);
INTERCONNECT SplitCLK_4_344_SplitCLK_2_343(net789_c1,net789);
INTERCONNECT SplitCLK_2_343_SplitCLK_6_339(net790_c1,net790);
INTERCONNECT SplitCLK_2_343_SplitCLK_4_342(net791_c1,net791);
INTERCONNECT SplitCLK_4_342_SplitCLK_4_340(net792_c1,net792);
INTERCONNECT SplitCLK_4_342_SplitCLK_2_341(net793_c1,net793);
INTERCONNECT SplitCLK_2_341_AND2T_38_n62(net794_c1,net794);
INTERCONNECT SplitCLK_2_341_DFFT_209__FPB_n602(net795_c1,net795);
INTERCONNECT SplitCLK_4_340_DFFT_210__FPB_n603(net796_c1,net796);
INTERCONNECT SplitCLK_4_340_DFFT_211__FPB_n604(net797_c1,net797);
INTERCONNECT SplitCLK_6_339_SplitCLK_4_337(net798_c1,net798);
INTERCONNECT SplitCLK_6_339_SplitCLK_4_338(net799_c1,net799);
INTERCONNECT SplitCLK_4_338_AND2T_14_n38(net800_c1,net800);
INTERCONNECT SplitCLK_4_338_OR2T_47_n71(net801_c1,net801);
INTERCONNECT SplitCLK_4_337_DFFT_161__FPB_n554(net802_c1,net802);
INTERCONNECT SplitCLK_4_337_DFFT_162__FPB_n555(net803_c1,net803);
INTERCONNECT SplitCLK_4_336_SplitCLK_6_332(net804_c1,net804);
INTERCONNECT SplitCLK_4_336_SplitCLK_4_335(net805_c1,net805);
INTERCONNECT SplitCLK_4_335_SplitCLK_4_333(net806_c1,net806);
INTERCONNECT SplitCLK_4_335_SplitCLK_4_334(net807_c1,net807);
INTERCONNECT SplitCLK_4_334_DFFT_160__FPB_n553(net808_c1,net808);
INTERCONNECT SplitCLK_4_334_DFFT_147__FPB_n540(net809_c1,net809);
INTERCONNECT SplitCLK_4_333_DFFT_212__FPB_n605(net810_c1,net810);
INTERCONNECT SplitCLK_4_333_DFFT_213__FPB_n606(net811_c1,net811);
INTERCONNECT SplitCLK_6_332_SplitCLK_4_330(net812_c1,net812);
INTERCONNECT SplitCLK_6_332_SplitCLK_0_331(net813_c1,net813);
INTERCONNECT SplitCLK_0_331_NOTT_18_n42(net814_c1,net814);
INTERCONNECT SplitCLK_0_331_DFFT_148__FPB_n541(net815_c1,net815);
INTERCONNECT SplitCLK_4_330_AND2T_12_n36(net816_c1,net816);
INTERCONNECT SplitCLK_4_330_AND2T_13_n37(net817_c1,net817);
INTERCONNECT SplitCLK_6_329_SplitCLK_0_321(net818_c1,net818);
INTERCONNECT SplitCLK_6_329_SplitCLK_2_328(net819_c1,net819);
INTERCONNECT SplitCLK_2_328_SplitCLK_2_324(net820_c1,net820);
INTERCONNECT SplitCLK_2_328_SplitCLK_4_327(net821_c1,net821);
INTERCONNECT SplitCLK_4_327_SplitCLK_4_325(net822_c1,net822);
INTERCONNECT SplitCLK_4_327_SplitCLK_4_326(net823_c1,net823);
INTERCONNECT SplitCLK_4_326_AND2T_55_n79(net824_c1,net824);
INTERCONNECT SplitCLK_4_326_OR2T_42_n66(net825_c1,net825);
INTERCONNECT SplitCLK_4_325_AND2T_16_n40(net826_c1,net826);
INTERCONNECT SplitCLK_4_325_AND2T_41_n65(net827_c1,net827);
INTERCONNECT SplitCLK_2_324_SplitCLK_4_322(net828_c1,net828);
INTERCONNECT SplitCLK_2_324_SplitCLK_4_323(net829_c1,net829);
INTERCONNECT SplitCLK_4_323_AND2T_80_n104(net830_c1,net830);
INTERCONNECT SplitCLK_4_323_AND2T_79_n103(net831_c1,net831);
INTERCONNECT SplitCLK_4_322_AND2T_56_n80(net832_c1,net832);
INTERCONNECT SplitCLK_4_322_OR2T_96_n120(net833_c1,net833);
INTERCONNECT SplitCLK_0_321_SplitCLK_6_317(net834_c1,net834);
INTERCONNECT SplitCLK_0_321_SplitCLK_4_320(net835_c1,net835);
INTERCONNECT SplitCLK_4_320_SplitCLK_4_318(net836_c1,net836);
INTERCONNECT SplitCLK_4_320_SplitCLK_4_319(net837_c1,net837);
INTERCONNECT SplitCLK_4_319_DFFT_150__FPB_n543(net838_c1,net838);
INTERCONNECT SplitCLK_4_319_DFFT_185__FPB_n578(net839_c1,net839);
INTERCONNECT SplitCLK_4_318_NOTT_11_n35(net840_c1,net840);
INTERCONNECT SplitCLK_4_318_DFFT_184__FPB_n577(net841_c1,net841);
INTERCONNECT SplitCLK_6_317_SplitCLK_4_315(net842_c1,net842);
INTERCONNECT SplitCLK_6_317_SplitCLK_4_316(net843_c1,net843);
INTERCONNECT SplitCLK_4_316_DFFT_163__FPB_n556(net844_c1,net844);
INTERCONNECT SplitCLK_4_316_DFFT_194__FPB_n587(net845_c1,net845);
INTERCONNECT SplitCLK_4_315_OR2T_75_n99(net846_c1,net846);
INTERCONNECT SplitCLK_4_315_DFFT_175__FPB_n568(net847_c1,net847);
INTERCONNECT SplitCLK_6_314_SplitCLK_0_283(net848_c1,net848);
INTERCONNECT SplitCLK_6_314_SplitCLK_2_313(net849_c1,net849);
INTERCONNECT SplitCLK_2_313_SplitCLK_6_298(net850_c1,net850);
INTERCONNECT SplitCLK_2_313_SplitCLK_4_312(net851_c1,net851);
INTERCONNECT SplitCLK_4_312_SplitCLK_0_305(net852_c1,net852);
INTERCONNECT SplitCLK_4_312_SplitCLK_2_311(net853_c1,net853);
INTERCONNECT SplitCLK_2_311_SplitCLK_2_308(net854_c1,net854);
INTERCONNECT SplitCLK_2_311_SplitCLK_4_310(net855_c1,net855);
INTERCONNECT SplitCLK_4_310_SplitCLK_2_503(net856_c1,net856);
INTERCONNECT SplitCLK_4_310_SplitCLK_4_309(net857_c1,net857);
INTERCONNECT SplitCLK_4_309_OR2T_111_n135(net858_c1,net858);
INTERCONNECT SplitCLK_4_309_DFFT_146__FPB_n539(net859_c1,net859);
INTERCONNECT SplitCLK_2_308_SplitCLK_4_306(net860_c1,net860);
INTERCONNECT SplitCLK_2_308_SplitCLK_4_307(net861_c1,net861);
INTERCONNECT SplitCLK_4_307_OR2T_100_n124(net862_c1,net862);
INTERCONNECT SplitCLK_4_307_DFFT_226__FPB_n619(net863_c1,net863);
INTERCONNECT SplitCLK_4_306_OR2T_112_n136(net864_c1,net864);
INTERCONNECT SplitCLK_4_306_DFFT_218__FPB_n611(net865_c1,net865);
INTERCONNECT SplitCLK_0_305_SplitCLK_4_301(net866_c1,net866);
INTERCONNECT SplitCLK_0_305_SplitCLK_4_304(net867_c1,net867);
INTERCONNECT SplitCLK_4_304_SplitCLK_4_302(net868_c1,net868);
INTERCONNECT SplitCLK_4_304_SplitCLK_4_303(net869_c1,net869);
INTERCONNECT SplitCLK_4_303_AND2T_110_n134(net870_c1,net870);
INTERCONNECT SplitCLK_4_303_OR2T_97_n121(net871_c1,net871);
INTERCONNECT SplitCLK_4_302_DFFT_220__FPB_n613(net872_c1,net872);
INTERCONNECT SplitCLK_4_302_DFFT_186__FPB_n579(net873_c1,net873);
INTERCONNECT SplitCLK_4_301_SplitCLK_4_299(net874_c1,net874);
INTERCONNECT SplitCLK_4_301_SplitCLK_4_300(net875_c1,net875);
INTERCONNECT SplitCLK_4_300_AND2T_101_n125(net876_c1,net876);
INTERCONNECT SplitCLK_4_300_OR2T_113_n137(net877_c1,net877);
INTERCONNECT SplitCLK_4_299_OR2T_93_n117(net878_c1,net878);
INTERCONNECT SplitCLK_4_299_DFFT_216__FPB_n609(net879_c1,net879);
INTERCONNECT SplitCLK_6_298_SplitCLK_0_290(net880_c1,net880);
INTERCONNECT SplitCLK_6_298_SplitCLK_2_297(net881_c1,net881);
INTERCONNECT SplitCLK_2_297_SplitCLK_6_293(net882_c1,net882);
INTERCONNECT SplitCLK_2_297_SplitCLK_4_296(net883_c1,net883);
INTERCONNECT SplitCLK_4_296_SplitCLK_4_294(net884_c1,net884);
INTERCONNECT SplitCLK_4_296_SplitCLK_4_295(net885_c1,net885);
INTERCONNECT SplitCLK_4_295_OR2T_104_n128(net886_c1,net886);
INTERCONNECT SplitCLK_4_295_DFFT_219__FPB_n612(net887_c1,net887);
INTERCONNECT SplitCLK_4_294_AND2T_103_n127(net888_c1,net888);
INTERCONNECT SplitCLK_4_294_AND2T_17_n41(net889_c1,net889);
INTERCONNECT SplitCLK_6_293_SplitCLK_4_291(net890_c1,net890);
INTERCONNECT SplitCLK_6_293_SplitCLK_4_292(net891_c1,net891);
INTERCONNECT SplitCLK_4_292_DFFT_254_state_obs2(net892_c1,net892);
INTERCONNECT SplitCLK_4_292_DFFT_253__FPB_n646(net893_c1,net893);
INTERCONNECT SplitCLK_4_291_DFFT_233__FPB_n626(net894_c1,net894);
INTERCONNECT SplitCLK_4_291_DFFT_252__FPB_n645(net895_c1,net895);
INTERCONNECT SplitCLK_0_290_SplitCLK_6_286(net896_c1,net896);
INTERCONNECT SplitCLK_0_290_SplitCLK_2_289(net897_c1,net897);
INTERCONNECT SplitCLK_2_289_SplitCLK_4_287(net898_c1,net898);
INTERCONNECT SplitCLK_2_289_SplitCLK_4_288(net899_c1,net899);
INTERCONNECT SplitCLK_4_288_OR2T_116_n140(net900_c1,net900);
INTERCONNECT SplitCLK_4_288_AND2T_98_n122(net901_c1,net901);
INTERCONNECT SplitCLK_4_287_AND2T_108_n132(net902_c1,net902);
INTERCONNECT SplitCLK_4_287_DFFT_217__FPB_n610(net903_c1,net903);
INTERCONNECT SplitCLK_6_286_SplitCLK_4_284(net904_c1,net904);
INTERCONNECT SplitCLK_6_286_SplitCLK_4_285(net905_c1,net905);
INTERCONNECT SplitCLK_4_285_DFFT_250__FPB_n643(net906_c1,net906);
INTERCONNECT SplitCLK_4_285_DFFT_251__FPB_n644(net907_c1,net907);
INTERCONNECT SplitCLK_4_284_NOTT_27_n51(net908_c1,net908);
INTERCONNECT SplitCLK_4_284_DFFT_249__FPB_n642(net909_c1,net909);
INTERCONNECT SplitCLK_0_283_SplitCLK_6_267(net910_c1,net910);
INTERCONNECT SplitCLK_0_283_SplitCLK_4_282(net911_c1,net911);
INTERCONNECT SplitCLK_4_282_SplitCLK_4_274(net912_c1,net912);
INTERCONNECT SplitCLK_4_282_SplitCLK_2_281(net913_c1,net913);
INTERCONNECT SplitCLK_2_281_SplitCLK_6_277(net914_c1,net914);
INTERCONNECT SplitCLK_2_281_SplitCLK_4_280(net915_c1,net915);
INTERCONNECT SplitCLK_4_280_SplitCLK_4_278(net916_c1,net916);
INTERCONNECT SplitCLK_4_280_SplitCLK_4_279(net917_c1,net917);
INTERCONNECT SplitCLK_4_279_DFFT_206__FPB_n599(net918_c1,net918);
INTERCONNECT SplitCLK_4_279_OR2T_76_n100(net919_c1,net919);
INTERCONNECT SplitCLK_4_278_AND2T_81_n105(net920_c1,net920);
INTERCONNECT SplitCLK_4_278_DFFT_201__FPB_n594(net921_c1,net921);
INTERCONNECT SplitCLK_6_277_SplitCLK_4_275(net922_c1,net922);
INTERCONNECT SplitCLK_6_277_SplitCLK_4_276(net923_c1,net923);
INTERCONNECT SplitCLK_4_276_AND2T_102_n126(net924_c1,net924);
INTERCONNECT SplitCLK_4_276_DFFT_200__FPB_n593(net925_c1,net925);
INTERCONNECT SplitCLK_4_275_DFFT_140__FBL_n533(net926_c1,net926);
INTERCONNECT SplitCLK_4_275_DFFT_135__FBL_n528(net927_c1,net927);
INTERCONNECT SplitCLK_4_274_SplitCLK_0_270(net928_c1,net928);
INTERCONNECT SplitCLK_4_274_SplitCLK_6_273(net929_c1,net929);
INTERCONNECT SplitCLK_6_273_SplitCLK_4_271(net930_c1,net930);
INTERCONNECT SplitCLK_6_273_SplitCLK_4_272(net931_c1,net931);
INTERCONNECT SplitCLK_4_272_DFFT_207__FPB_n600(net932_c1,net932);
INTERCONNECT SplitCLK_4_272_DFFT_196__FPB_n589(net933_c1,net933);
INTERCONNECT SplitCLK_4_271_AND2T_77_n101(net934_c1,net934);
INTERCONNECT SplitCLK_4_271_OR2T_94_n118(net935_c1,net935);
INTERCONNECT SplitCLK_0_270_SplitCLK_4_268(net936_c1,net936);
INTERCONNECT SplitCLK_0_270_SplitCLK_0_269(net937_c1,net937);
INTERCONNECT SplitCLK_0_269_DFFT_199__FPB_n592(net938_c1,net938);
INTERCONNECT SplitCLK_0_269_DFFT_198__FPB_n591(net939_c1,net939);
INTERCONNECT SplitCLK_4_268_AND2T_78_n102(net940_c1,net940);
INTERCONNECT SplitCLK_4_268_AND2T_95_n119(net941_c1,net941);
INTERCONNECT SplitCLK_6_267_SplitCLK_4_259(net942_c1,net942);
INTERCONNECT SplitCLK_6_267_SplitCLK_2_266(net943_c1,net943);
INTERCONNECT SplitCLK_2_266_SplitCLK_6_262(net944_c1,net944);
INTERCONNECT SplitCLK_2_266_SplitCLK_4_265(net945_c1,net945);
INTERCONNECT SplitCLK_4_265_SplitCLK_4_263(net946_c1,net946);
INTERCONNECT SplitCLK_4_265_SplitCLK_4_264(net947_c1,net947);
INTERCONNECT SplitCLK_4_264_AND2T_107_n131(net948_c1,net948);
INTERCONNECT SplitCLK_4_264_DFFT_215__FPB_n608(net949_c1,net949);
INTERCONNECT SplitCLK_4_263_DFFT_214__FPB_n607(net950_c1,net950);
INTERCONNECT SplitCLK_4_263_DFFT_144__FBL_n537(net951_c1,net951);
INTERCONNECT SplitCLK_6_262_SplitCLK_4_260(net952_c1,net952);
INTERCONNECT SplitCLK_6_262_SplitCLK_4_261(net953_c1,net953);
INTERCONNECT SplitCLK_4_261_DFFT_259_state_obs3(net954_c1,net954);
INTERCONNECT SplitCLK_4_261_OR2T_106_n130(net955_c1,net955);
INTERCONNECT SplitCLK_4_260_DFFT_255__FPB_n648(net956_c1,net956);
INTERCONNECT SplitCLK_4_260_DFFT_258__FPB_n651(net957_c1,net957);
INTERCONNECT SplitCLK_4_259_SplitCLK_4_255(net958_c1,net958);
INTERCONNECT SplitCLK_4_259_SplitCLK_0_258(net959_c1,net959);
INTERCONNECT SplitCLK_0_258_SplitCLK_4_256(net960_c1,net960);
INTERCONNECT SplitCLK_0_258_SplitCLK_0_257(net961_c1,net961);
INTERCONNECT SplitCLK_0_257_DFFT_132__PIPL_n183(net962_c1,net962);
INTERCONNECT SplitCLK_0_257_DFFT_223__FPB_n616(net963_c1,net963);
INTERCONNECT SplitCLK_4_256_OR2T_105_n129(net964_c1,net964);
INTERCONNECT SplitCLK_4_256_DFFT_197__FPB_n590(net965_c1,net965);
INTERCONNECT SplitCLK_4_255_SplitCLK_4_253(net966_c1,net966);
INTERCONNECT SplitCLK_4_255_SplitCLK_4_254(net967_c1,net967);
INTERCONNECT SplitCLK_4_254_NOTT_115_n139(net968_c1,net968);
INTERCONNECT SplitCLK_4_254_DFFT_257__FPB_n650(net969_c1,net969);
INTERCONNECT SplitCLK_4_253_DFFT_131__PIPL_n182(net970_c1,net970);
INTERCONNECT SplitCLK_4_253_DFFT_256__FPB_n649(net971_c1,net971);
INTERCONNECT GCLK_Pad_SplitCLK_0_507(GCLK_Pad,net972);
INTERCONNECT Split_HOLD_621_DFFT_217__FPB_n610(net973_c1,net973);
INTERCONNECT Split_HOLD_622_DFFT_223__FPB_n616(net974_c1,net974);

endmodule
