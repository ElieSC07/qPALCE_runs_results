module TAP_route(
input GCLK_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output state_obs2_Pad,
output state_obs3_Pad);

wire net0_c1;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire TRST_Pad;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire state_obs0_Pad;
wire net136_c1;
wire state_obs1_Pad;
wire net137_c1;
wire state_obs2_Pad;
wire net138_c1;
wire state_obs3_Pad;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire GCLK_Pad;
wire net353;

XOR2T XOR2T_28_n52(net229,net4,net23,net11_c1);
DFFT DFFT_83_state_obs1(net249,net130,net136_c1);
DFFT DFFT_91_state_obs3(net331,net129,net138_c1);
NOTT NOTT_8_n32(net188,net86,net1_c1);
NOTT NOTT_9_n33(net187,net68,net3_c1);
DFFT DFFT_39_state0_buf(net186,net90,net139_c1);
AND2T AND2T_20_n44(net201,net8,net17,net12_c1);
AND2T AND2T_12_n36(net185,net75,net104,net13_c1);
AND2T AND2T_23_n47(net209,net16,net103,net23_c1);
AND2T AND2T_32_n56(net184,net22,net123,net25_c1);
AND2T AND2T_33_n57(net341,net25,net126,net27_c1);
AND2T AND2T_25_n49(net183,net35,net107,net28_c1);
AND2T AND2T_26_n50(net182,net28,net26,net4_c1);
AND2T AND2T_27_n51(net225,net11,net117,net7_c1);
AND2T AND2T_19_n43(net283,net5,net101,net8_c1);
AND2T AND2T_36_n60(net181,net82,net110,net10_c1);
AND2T AND2T_37_n61(net284,net10,net30,net14_c1);
AND2T AND2T_29_n53(net180,net81,net71,net15_c1);
AND2T AND2T_38_n62(net179,net14,net29,net18_c1);
DFFT DFFT_79_state_obs0(net178,net120,net135_c1);
DFFT DFFT_87_state_obs2(net269,net119,net137_c1);
OR2T OR2T_11_n35(net230,net72,net66,net9_c1);
OR2T OR2T_21_n45(net177,net61,net64,net16_c1);
OR2T OR2T_13_n37(net176,net13,net114,net17_c1);
OR2T OR2T_30_n54(net259,net15,net121,net19_c1);
OR2T OR2T_22_n46(net210,net49,net39,net20_c1);
OR2T OR2T_31_n55(net323,net63,net69,net22_c1);
OR2T OR2T_15_n39(net175,net36,net118,net24_c1);
OR2T OR2T_24_n48(net174,net31,net42,net26_c1);
OR2T OR2T_17_n41(net311,net65,net122,net2_c1);
OR2T OR2T_18_n42(net307,net2,net24,net5_c1);
OR2T OR2T_34_n58(net219,net45,net102,net29_c1);
OR2T OR2T_35_n59(net291,net70,net106,net30_c1);
DFFT DFFT_47__ADJFBL_n194(net173,net67,net90_c1);
DFFT DFFT_40_state1_buf(net172,net91,net140_c1);
NOTT NOTT_10_n34(net171,net77,net6_c1);
NOTT NOTT_14_n38(net170,net60,net21_c1);
NOTT NOTT_16_n40(net169,net85,net0_c1);
DFFT DFFT_48__ADJFBL_n195(net168,net73,net91_c1);
DFFT DFFT_41_state2_buf(net332,net92,net141_c1);
DFFT DFFT_49__ADJFBL_n196(net167,net97,net92_c1);
DFFT DFFT_42_state3_buf(net166,net55,net142_c1);
DFFT DFFT_50__FBL_n197(net220,net99,net94_c1);
DFFT DFFT_51__FBL_n198(net165,net37,net95_c1);
DFFT DFFT_52__FBL_n199(net241,net44,net96_c1);
DFFT DFFT_60__FPB_n207(net164,net109,net114_c1);
DFFT DFFT_43__PIPL_n76(net242,net139,net131_c1);
DFFT DFFT_53__FBL_n200(net324,net100,net93_c1);
DFFT DFFT_61__FPB_n208(net226,net52,net118_c1);
DFFT DFFT_44__PIPL_n77(net265,net140,net132_c1);
DFFT DFFT_54__FPB_n201(net342,net76,net97_c1);
DFFT DFFT_70__FPB_n217(net163,net89,net121_c1);
DFFT DFFT_62__FPB_n209(net308,net57,net122_c1);
DFFT DFFT_45__PIPL_n78(net162,net141,net133_c1);
DFFT DFFT_63__FPB_n210(net161,net51,net98_c1);
DFFT DFFT_55__FPB_n202(net160,net18,net99_c1);
DFFT DFFT_71__FPB_n218(net301,net54,net123_c1);
DFFT DFFT_46__PIPL_n79(net347,net142,net134_c1);
DFFT DFFT_64__FPB_n211(net159,net98,net101_c1);
DFFT DFFT_56__FPB_n203(net158,net48,net100_c1);
DFFT DFFT_80__FPB_n227(net157,net132,net125_c1);
DFFT DFFT_72__FPB_n219(net156,net19,net126_c1);
DFFT DFFT_73__FPB_n220(net155,net32,net102_c1);
DFFT DFFT_65__FPB_n212(net154,net40,net103_c1);
DFFT DFFT_57__FPB_n204(net153,net62,net104_c1);
DFFT DFFT_81__FPB_n228(net152,net125,net128_c1);
DFFT DFFT_74__FPB_n221(net292,net59,net106_c1);
DFFT DFFT_66__FPB_n213(net260,net41,net107_c1);
DFFT DFFT_58__FPB_n205(net202,net87,net105_c1);
DFFT DFFT_90__FPB_n237(net351,net127,net129_c1);
DFFT DFFT_82__FPB_n229(net266,net128,net130_c1);
SPLITT Split_100_n247(net21,net46_c1,net78_c1);
SPLITT Split_101_n248(net78,net51_c1,net82_c1);
SPLITT Split_102_n249(net46,net54_c1,net84_c1);
SPLITT Split_110_n257(net80,net55_c1,net85_c1);
SPLITT Split_103_n250(net0,net33_c1,net63_c1);
SPLITT Split_111_n258(net50,net56_c1,net87_c1);
SPLITT Split_104_n251(net33,net35_c1,net65_c1);
SPLITT Split_112_n259(net95,net58_c1,net88_c1);
SPLITT Split_120_n267(net53,net59_c1,net89_c1);
SPLITT Split_105_n252(net12,net37_c1,net67_c1);
SPLITT Split_113_n260(net88,net39_c1,net68_c1);
SPLITT Split_106_n253(net20,net40_c1,net70_c1);
SPLITT Split_114_n261(net58,net41_c1,net71_c1);
SPLITT Split_107_n254(net7,net44_c1,net73_c1);
SPLITT Split_115_n262(net96,net43_c1,net74_c1);
SPLITT Split_108_n255(net27,net48_c1,net76_c1);
SPLITT Split_116_n263(net74,net49_c1,net77_c1);
SPLITT Split_109_n256(net94,net50_c1,net80_c1);
SPLITT Split_117_n264(net43,net52_c1,net81_c1);
SPLITT Split_118_n265(net93,net53_c1,net83_c1);
SPLITT Split_119_n266(net83,net57_c1,net86_c1);
DFFT DFFT_75__FPB_n222(net151,net56,net110_c1);
DFFT DFFT_67__FPB_n214(net150,net84,net108_c1);
DFFT DFFT_59__FPB_n206(net149,net105,net109_c1);
DFFT DFFT_84__FPB_n231(net148,net133,net111_c1);
DFFT DFFT_76__FPB_n223(net147,net131,net112_c1);
DFFT DFFT_68__FPB_n215(net302,net108,net113_c1);
DFFT DFFT_85__FPB_n232(net270,net111,net115_c1);
DFFT DFFT_77__FPB_n224(net250,net112,net116_c1);
DFFT DFFT_69__FPB_n216(net312,net113,net117_c1);
DFFT DFFT_86__FPB_n233(net146,net115,net119_c1);
DFFT DFFT_78__FPB_n225(net145,net116,net120_c1);
SPLITT Split_92_n239(net1,net47_c1,net79_c1);
SPLITT Split_93_n240(net79,net31_c1,net61_c1);
SPLITT Split_94_n241(net47,net32_c1,net62_c1);
SPLITT Split_95_n242(net3,net34_c1,net64_c1);
SPLITT Split_96_n243(net34,net36_c1,net66_c1);
SPLITT Split_97_n244(net6,net38_c1,net69_c1);
SPLITT Split_98_n245(net38,net42_c1,net72_c1);
SPLITT Split_99_n246(net9,net45_c1,net75_c1);
DFFT DFFT_88__FPB_n235(net348,net134,net124_c1);
DFFT DFFT_89__FPB_n236(net352,net124,net127_c1);
SPLITT SplitCLK_4_85(net350,net352_c1,net351_c1);
SPLITT SplitCLK_4_86(net343,net350_c1,net349_c1);
SPLITT SplitCLK_4_87(net346,net348_c1,net347_c1);
SPLITT SplitCLK_6_88(net344,net346_c1,net345_c1);
SPLITT SplitCLK_4_89(net333,net344_c1,net343_c1);
SPLITT SplitCLK_4_90(net340,net342_c1,net341_c1);
SPLITT SplitCLK_0_91(net335,net340_c1,net339_c1);
SPLITT SplitCLK_4_92(net336,net337_c1,net338_c1);
SPLITT SplitCLK_4_93(net334,net336_c1,net335_c1);
SPLITT SplitCLK_6_94(net313,net333_c1,net334_c1);
SPLITT SplitCLK_4_95(net330,net331_c1,net332_c1);
SPLITT SplitCLK_2_96(net325,net329_c1,net330_c1);
SPLITT SplitCLK_6_97(net326,net327_c1,net328_c1);
SPLITT SplitCLK_6_98(net315,net325_c1,net326_c1);
SPLITT SplitCLK_4_99(net322,net323_c1,net324_c1);
SPLITT SplitCLK_4_100(net317,net321_c1,net322_c1);
SPLITT SplitCLK_6_101(net318,net320_c1,net319_c1);
SPLITT SplitCLK_4_102(net316,net318_c1,net317_c1);
SPLITT SplitCLK_6_103(net314,net316_c1,net315_c1);
SPLITT SplitCLK_6_104(net271,net313_c1,net314_c1);
SPLITT SplitCLK_4_105(net310,net311_c1,net312_c1);
SPLITT SplitCLK_4_106(net303,net310_c1,net309_c1);
SPLITT SplitCLK_4_107(net306,net308_c1,net307_c1);
SPLITT SplitCLK_2_108(net304,net305_c1,net306_c1);
SPLITT SplitCLK_4_109(net293,net304_c1,net303_c1);
SPLITT SplitCLK_4_110(net300,net301_c1,net302_c1);
SPLITT SplitCLK_0_111(net295,net300_c1,net299_c1);
SPLITT SplitCLK_4_112(net296,net297_c1,net298_c1);
SPLITT SplitCLK_4_113(net294,net296_c1,net295_c1);
SPLITT SplitCLK_0_114(net273,net293_c1,net294_c1);
SPLITT SplitCLK_4_115(net290,net291_c1,net292_c1);
SPLITT SplitCLK_0_116(net285,net290_c1,net289_c1);
SPLITT SplitCLK_6_117(net286,net287_c1,net288_c1);
SPLITT SplitCLK_6_118(net275,net285_c1,net286_c1);
SPLITT SplitCLK_4_119(net282,net284_c1,net283_c1);
SPLITT SplitCLK_4_120(net277,net282_c1,net281_c1);
SPLITT SplitCLK_2_121(net278,net280_c1,net279_c1);
SPLITT SplitCLK_4_122(net276,net278_c1,net277_c1);
SPLITT SplitCLK_2_123(net274,net276_c1,net275_c1);
SPLITT SplitCLK_4_124(net272,net274_c1,net273_c1);
SPLITT SplitCLK_0_125(net143,net271_c1,net272_c1);
SPLITT SplitCLK_0_126(net268,net269_c1,net270_c1);
SPLITT SplitCLK_0_127(net261,net268_c1,net267_c1);
SPLITT SplitCLK_4_128(net264,net266_c1,net265_c1);
SPLITT SplitCLK_2_129(net262,net263_c1,net264_c1);
SPLITT SplitCLK_6_130(net251,net261_c1,net262_c1);
SPLITT SplitCLK_4_131(net258,net260_c1,net259_c1);
SPLITT SplitCLK_4_132(net253,net257_c1,net258_c1);
SPLITT SplitCLK_2_133(net254,net255_c1,net256_c1);
SPLITT SplitCLK_0_134(net252,net254_c1,net253_c1);
SPLITT SplitCLK_4_135(net231,net251_c1,net252_c1);
SPLITT SplitCLK_4_136(net248,net250_c1,net249_c1);
SPLITT SplitCLK_0_137(net243,net248_c1,net247_c1);
SPLITT SplitCLK_6_138(net244,net246_c1,net245_c1);
SPLITT SplitCLK_6_139(net233,net243_c1,net244_c1);
SPLITT SplitCLK_4_140(net240,net242_c1,net241_c1);
SPLITT SplitCLK_4_141(net235,net240_c1,net239_c1);
SPLITT SplitCLK_6_142(net236,net237_c1,net238_c1);
SPLITT SplitCLK_4_143(net234,net236_c1,net235_c1);
SPLITT SplitCLK_6_144(net232,net233_c1,net234_c1);
SPLITT SplitCLK_6_145(net189,net231_c1,net232_c1);
SPLITT SplitCLK_4_146(net228,net229_c1,net230_c1);
SPLITT SplitCLK_2_147(net221,net227_c1,net228_c1);
SPLITT SplitCLK_0_148(net224,net225_c1,net226_c1);
SPLITT SplitCLK_2_149(net222,net223_c1,net224_c1);
SPLITT SplitCLK_4_150(net211,net222_c1,net221_c1);
SPLITT SplitCLK_4_151(net218,net220_c1,net219_c1);
SPLITT SplitCLK_0_152(net213,net218_c1,net217_c1);
SPLITT SplitCLK_4_153(net214,net215_c1,net216_c1);
SPLITT SplitCLK_4_154(net212,net214_c1,net213_c1);
SPLITT SplitCLK_0_155(net191,net211_c1,net212_c1);
SPLITT SplitCLK_4_156(net208,net209_c1,net210_c1);
SPLITT SplitCLK_4_157(net203,net208_c1,net207_c1);
SPLITT SplitCLK_6_158(net204,net205_c1,net206_c1);
SPLITT SplitCLK_6_159(net193,net203_c1,net204_c1);
SPLITT SplitCLK_4_160(net200,net201_c1,net202_c1);
SPLITT SplitCLK_2_161(net195,net199_c1,net200_c1);
SPLITT SplitCLK_6_162(net196,net197_c1,net198_c1);
SPLITT SplitCLK_4_163(net194,net196_c1,net195_c1);
SPLITT SplitCLK_2_164(net192,net194_c1,net193_c1);
SPLITT SplitCLK_4_165(net190,net192_c1,net191_c1);
SPLITT SplitCLK_2_166(net144,net190_c1,net189_c1);
wire dummy0;
SPLITT SplitCLK_2_167(net305,net188_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_2_168(net205,net187_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_4_169(net247,net186_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_4_170(net207,net185_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_171(net337,net184_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_4_172(net287,net183_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_2_173(net288,net182_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_4_174(net281,net181_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_2_175(net257,net180_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_4_176(net217,net179_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_2_177(net245,net178_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_2_178(net223,net177_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_2_179(net197,net176_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_2_180(net227,net175_c1,dummy13);
wire dummy14;
SPLITT SplitCLK_4_181(net289,net174_c1,dummy14);
wire dummy15;
SPLITT SplitCLK_4_182(net237,net173_c1,dummy15);
wire dummy16;
SPLITT SplitCLK_4_183(net267,net172_c1,dummy16);
wire dummy17;
SPLITT SplitCLK_4_184(net321,net171_c1,dummy17);
wire dummy18;
SPLITT SplitCLK_4_185(net299,net170_c1,dummy18);
wire dummy19;
SPLITT SplitCLK_4_186(net339,net169_c1,dummy19);
wire dummy20;
SPLITT SplitCLK_4_187(net255,net168_c1,dummy20);
wire dummy21;
SPLITT SplitCLK_2_188(net345,net167_c1,dummy21);
wire dummy22;
SPLITT SplitCLK_4_189(net349,net166_c1,dummy22);
wire dummy23;
SPLITT SplitCLK_4_190(net239,net165_c1,dummy23);
wire dummy24;
SPLITT SplitCLK_4_191(net198,net164_c1,dummy24);
wire dummy25;
SPLITT SplitCLK_2_192(net319,net163_c1,dummy25);
wire dummy26;
SPLITT SplitCLK_4_193(net327,net162_c1,dummy26);
wire dummy27;
SPLITT SplitCLK_2_194(net297,net161_c1,dummy27);
wire dummy28;
SPLITT SplitCLK_2_195(net215,net160_c1,dummy28);
wire dummy29;
SPLITT SplitCLK_2_196(net298,net159_c1,dummy29);
wire dummy30;
SPLITT SplitCLK_2_197(net338,net158_c1,dummy30);
wire dummy31;
SPLITT SplitCLK_2_198(net263,net157_c1,dummy31);
wire dummy32;
SPLITT SplitCLK_4_199(net320,net156_c1,dummy32);
wire dummy33;
SPLITT SplitCLK_2_200(net279,net155_c1,dummy33);
wire dummy34;
SPLITT SplitCLK_4_201(net206,net154_c1,dummy34);
wire dummy35;
SPLITT SplitCLK_2_202(net216,net153_c1,dummy35);
wire dummy36;
SPLITT SplitCLK_2_203(net256,net152_c1,dummy36);
wire dummy37;
SPLITT SplitCLK_4_204(net280,net151_c1,dummy37);
wire dummy38;
SPLITT SplitCLK_4_205(net309,net150_c1,dummy38);
wire dummy39;
SPLITT SplitCLK_2_206(net199,net149_c1,dummy39);
wire dummy40;
SPLITT SplitCLK_2_207(net329,net148_c1,dummy40);
wire dummy41;
SPLITT SplitCLK_2_208(net238,net147_c1,dummy41);
wire dummy42;
SPLITT SplitCLK_2_209(net328,net146_c1,dummy42);
wire dummy43;
SPLITT SplitCLK_4_210(net246,net145_c1,dummy43);
SPLITT SplitCLK_0_211(net353,net143_c1,net144_c1);
INTERCONNECT NOTT_16_n40_Split_103_n250(net0_c1,net0);
INTERCONNECT NOTT_8_n32_Split_92_n239(net1_c1,net1);
INTERCONNECT OR2T_17_n41_OR2T_18_n42(net2_c1,net2);
INTERCONNECT NOTT_9_n33_Split_95_n242(net3_c1,net3);
INTERCONNECT AND2T_26_n50_XOR2T_28_n52(net4_c1,net4);
INTERCONNECT OR2T_18_n42_AND2T_19_n43(net5_c1,net5);
INTERCONNECT NOTT_10_n34_Split_97_n244(net6_c1,net6);
INTERCONNECT AND2T_27_n51_Split_107_n254(net7_c1,net7);
INTERCONNECT AND2T_19_n43_AND2T_20_n44(net8_c1,net8);
INTERCONNECT OR2T_11_n35_Split_99_n246(net9_c1,net9);
INTERCONNECT AND2T_36_n60_AND2T_37_n61(net10_c1,net10);
INTERCONNECT XOR2T_28_n52_AND2T_27_n51(net11_c1,net11);
INTERCONNECT AND2T_20_n44_Split_105_n252(net12_c1,net12);
INTERCONNECT AND2T_12_n36_OR2T_13_n37(net13_c1,net13);
INTERCONNECT AND2T_37_n61_AND2T_38_n62(net14_c1,net14);
INTERCONNECT AND2T_29_n53_OR2T_30_n54(net15_c1,net15);
INTERCONNECT OR2T_21_n45_AND2T_23_n47(net16_c1,net16);
INTERCONNECT OR2T_13_n37_AND2T_20_n44(net17_c1,net17);
INTERCONNECT AND2T_38_n62_DFFT_55__FPB_n202(net18_c1,net18);
INTERCONNECT OR2T_30_n54_DFFT_72__FPB_n219(net19_c1,net19);
INTERCONNECT OR2T_22_n46_Split_106_n253(net20_c1,net20);
INTERCONNECT NOTT_14_n38_Split_100_n247(net21_c1,net21);
INTERCONNECT OR2T_31_n55_AND2T_32_n56(net22_c1,net22);
INTERCONNECT AND2T_23_n47_XOR2T_28_n52(net23_c1,net23);
INTERCONNECT OR2T_15_n39_OR2T_18_n42(net24_c1,net24);
INTERCONNECT AND2T_32_n56_AND2T_33_n57(net25_c1,net25);
INTERCONNECT OR2T_24_n48_AND2T_26_n50(net26_c1,net26);
INTERCONNECT AND2T_33_n57_Split_108_n255(net27_c1,net27);
INTERCONNECT AND2T_25_n49_AND2T_26_n50(net28_c1,net28);
INTERCONNECT OR2T_34_n58_AND2T_38_n62(net29_c1,net29);
INTERCONNECT OR2T_35_n59_AND2T_37_n61(net30_c1,net30);
INTERCONNECT Split_93_n240_OR2T_24_n48(net31_c1,net31);
INTERCONNECT Split_94_n241_DFFT_73__FPB_n220(net32_c1,net32);
INTERCONNECT Split_103_n250_Split_104_n251(net33_c1,net33);
INTERCONNECT Split_95_n242_Split_96_n243(net34_c1,net34);
INTERCONNECT Split_104_n251_AND2T_25_n49(net35_c1,net35);
INTERCONNECT Split_96_n243_OR2T_15_n39(net36_c1,net36);
INTERCONNECT Split_105_n252_DFFT_51__FBL_n198(net37_c1,net37);
INTERCONNECT Split_97_n244_Split_98_n245(net38_c1,net38);
INTERCONNECT Split_113_n260_OR2T_22_n46(net39_c1,net39);
INTERCONNECT Split_106_n253_DFFT_65__FPB_n212(net40_c1,net40);
INTERCONNECT Split_114_n261_DFFT_66__FPB_n213(net41_c1,net41);
INTERCONNECT Split_98_n245_OR2T_24_n48(net42_c1,net42);
INTERCONNECT Split_115_n262_Split_117_n264(net43_c1,net43);
INTERCONNECT Split_107_n254_DFFT_52__FBL_n199(net44_c1,net44);
INTERCONNECT Split_99_n246_OR2T_34_n58(net45_c1,net45);
INTERCONNECT Split_100_n247_Split_102_n249(net46_c1,net46);
INTERCONNECT Split_92_n239_Split_94_n241(net47_c1,net47);
INTERCONNECT Split_108_n255_DFFT_56__FPB_n203(net48_c1,net48);
INTERCONNECT Split_116_n263_OR2T_22_n46(net49_c1,net49);
INTERCONNECT Split_109_n256_Split_111_n258(net50_c1,net50);
INTERCONNECT Split_101_n248_DFFT_63__FPB_n210(net51_c1,net51);
INTERCONNECT Split_117_n264_DFFT_61__FPB_n208(net52_c1,net52);
INTERCONNECT Split_118_n265_Split_120_n267(net53_c1,net53);
INTERCONNECT Split_102_n249_DFFT_71__FPB_n218(net54_c1,net54);
INTERCONNECT Split_110_n257_DFFT_42_state3_buf(net55_c1,net55);
INTERCONNECT Split_111_n258_DFFT_75__FPB_n222(net56_c1,net56);
INTERCONNECT Split_119_n266_DFFT_62__FPB_n209(net57_c1,net57);
INTERCONNECT Split_112_n259_Split_114_n261(net58_c1,net58);
INTERCONNECT Split_120_n267_DFFT_74__FPB_n221(net59_c1,net59);
INTERCONNECT TRST_Pad_NOTT_14_n38(TRST_Pad,net60);
INTERCONNECT Split_93_n240_OR2T_21_n45(net61_c1,net61);
INTERCONNECT Split_94_n241_DFFT_57__FPB_n204(net62_c1,net62);
INTERCONNECT Split_103_n250_OR2T_31_n55(net63_c1,net63);
INTERCONNECT Split_95_n242_OR2T_21_n45(net64_c1,net64);
INTERCONNECT Split_104_n251_OR2T_17_n41(net65_c1,net65);
INTERCONNECT Split_96_n243_OR2T_11_n35(net66_c1,net66);
INTERCONNECT Split_105_n252_DFFT_47__ADJFBL_n194(net67_c1,net67);
INTERCONNECT Split_113_n260_NOTT_9_n33(net68_c1,net68);
INTERCONNECT Split_97_n244_OR2T_31_n55(net69_c1,net69);
INTERCONNECT Split_106_n253_OR2T_35_n59(net70_c1,net70);
INTERCONNECT Split_114_n261_AND2T_29_n53(net71_c1,net71);
INTERCONNECT Split_98_n245_OR2T_11_n35(net72_c1,net72);
INTERCONNECT Split_107_n254_DFFT_48__ADJFBL_n195(net73_c1,net73);
INTERCONNECT Split_115_n262_Split_116_n263(net74_c1,net74);
INTERCONNECT Split_99_n246_AND2T_12_n36(net75_c1,net75);
INTERCONNECT Split_108_n255_DFFT_54__FPB_n201(net76_c1,net76);
INTERCONNECT Split_116_n263_NOTT_10_n34(net77_c1,net77);
INTERCONNECT Split_100_n247_Split_101_n248(net78_c1,net78);
INTERCONNECT Split_92_n239_Split_93_n240(net79_c1,net79);
INTERCONNECT Split_109_n256_Split_110_n257(net80_c1,net80);
INTERCONNECT Split_117_n264_AND2T_29_n53(net81_c1,net81);
INTERCONNECT Split_101_n248_AND2T_36_n60(net82_c1,net82);
INTERCONNECT Split_118_n265_Split_119_n266(net83_c1,net83);
INTERCONNECT Split_102_n249_DFFT_67__FPB_n214(net84_c1,net84);
INTERCONNECT Split_110_n257_NOTT_16_n40(net85_c1,net85);
INTERCONNECT Split_119_n266_NOTT_8_n32(net86_c1,net86);
INTERCONNECT Split_111_n258_DFFT_58__FPB_n205(net87_c1,net87);
INTERCONNECT Split_112_n259_Split_113_n260(net88_c1,net88);
INTERCONNECT Split_120_n267_DFFT_70__FPB_n217(net89_c1,net89);
INTERCONNECT DFFT_47__ADJFBL_n194_DFFT_39_state0_buf(net90_c1,net90);
INTERCONNECT DFFT_48__ADJFBL_n195_DFFT_40_state1_buf(net91_c1,net91);
INTERCONNECT DFFT_49__ADJFBL_n196_DFFT_41_state2_buf(net92_c1,net92);
INTERCONNECT DFFT_53__FBL_n200_Split_118_n265(net93_c1,net93);
INTERCONNECT DFFT_50__FBL_n197_Split_109_n256(net94_c1,net94);
INTERCONNECT DFFT_51__FBL_n198_Split_112_n259(net95_c1,net95);
INTERCONNECT DFFT_52__FBL_n199_Split_115_n262(net96_c1,net96);
INTERCONNECT DFFT_54__FPB_n201_DFFT_49__ADJFBL_n196(net97_c1,net97);
INTERCONNECT DFFT_63__FPB_n210_DFFT_64__FPB_n211(net98_c1,net98);
INTERCONNECT DFFT_55__FPB_n202_DFFT_50__FBL_n197(net99_c1,net99);
INTERCONNECT DFFT_56__FPB_n203_DFFT_53__FBL_n200(net100_c1,net100);
INTERCONNECT DFFT_64__FPB_n211_AND2T_19_n43(net101_c1,net101);
INTERCONNECT DFFT_73__FPB_n220_OR2T_34_n58(net102_c1,net102);
INTERCONNECT DFFT_65__FPB_n212_AND2T_23_n47(net103_c1,net103);
INTERCONNECT DFFT_57__FPB_n204_AND2T_12_n36(net104_c1,net104);
INTERCONNECT DFFT_58__FPB_n205_DFFT_59__FPB_n206(net105_c1,net105);
INTERCONNECT DFFT_74__FPB_n221_OR2T_35_n59(net106_c1,net106);
INTERCONNECT DFFT_66__FPB_n213_AND2T_25_n49(net107_c1,net107);
INTERCONNECT DFFT_67__FPB_n214_DFFT_68__FPB_n215(net108_c1,net108);
INTERCONNECT DFFT_59__FPB_n206_DFFT_60__FPB_n207(net109_c1,net109);
INTERCONNECT DFFT_75__FPB_n222_AND2T_36_n60(net110_c1,net110);
INTERCONNECT DFFT_84__FPB_n231_DFFT_85__FPB_n232(net111_c1,net111);
INTERCONNECT DFFT_76__FPB_n223_DFFT_77__FPB_n224(net112_c1,net112);
INTERCONNECT DFFT_68__FPB_n215_DFFT_69__FPB_n216(net113_c1,net113);
INTERCONNECT DFFT_60__FPB_n207_OR2T_13_n37(net114_c1,net114);
INTERCONNECT DFFT_85__FPB_n232_DFFT_86__FPB_n233(net115_c1,net115);
INTERCONNECT DFFT_77__FPB_n224_DFFT_78__FPB_n225(net116_c1,net116);
INTERCONNECT DFFT_69__FPB_n216_AND2T_27_n51(net117_c1,net117);
INTERCONNECT DFFT_61__FPB_n208_OR2T_15_n39(net118_c1,net118);
INTERCONNECT DFFT_86__FPB_n233_DFFT_87_state_obs2(net119_c1,net119);
INTERCONNECT DFFT_78__FPB_n225_DFFT_79_state_obs0(net120_c1,net120);
INTERCONNECT DFFT_70__FPB_n217_OR2T_30_n54(net121_c1,net121);
INTERCONNECT DFFT_62__FPB_n209_OR2T_17_n41(net122_c1,net122);
INTERCONNECT DFFT_71__FPB_n218_AND2T_32_n56(net123_c1,net123);
INTERCONNECT DFFT_88__FPB_n235_DFFT_89__FPB_n236(net124_c1,net124);
INTERCONNECT DFFT_80__FPB_n227_DFFT_81__FPB_n228(net125_c1,net125);
INTERCONNECT DFFT_72__FPB_n219_AND2T_33_n57(net126_c1,net126);
INTERCONNECT DFFT_89__FPB_n236_DFFT_90__FPB_n237(net127_c1,net127);
INTERCONNECT DFFT_81__FPB_n228_DFFT_82__FPB_n229(net128_c1,net128);
INTERCONNECT DFFT_90__FPB_n237_DFFT_91_state_obs3(net129_c1,net129);
INTERCONNECT DFFT_82__FPB_n229_DFFT_83_state_obs1(net130_c1,net130);
INTERCONNECT DFFT_43__PIPL_n76_DFFT_76__FPB_n223(net131_c1,net131);
INTERCONNECT DFFT_44__PIPL_n77_DFFT_80__FPB_n227(net132_c1,net132);
INTERCONNECT DFFT_45__PIPL_n78_DFFT_84__FPB_n231(net133_c1,net133);
INTERCONNECT DFFT_46__PIPL_n79_DFFT_88__FPB_n235(net134_c1,net134);
INTERCONNECT DFFT_79_state_obs0_state_obs0_Pad(net135_c1,state_obs0_Pad);
INTERCONNECT DFFT_83_state_obs1_state_obs1_Pad(net136_c1,state_obs1_Pad);
INTERCONNECT DFFT_87_state_obs2_state_obs2_Pad(net137_c1,state_obs2_Pad);
INTERCONNECT DFFT_91_state_obs3_state_obs3_Pad(net138_c1,state_obs3_Pad);
INTERCONNECT DFFT_39_state0_buf_DFFT_43__PIPL_n76(net139_c1,net139);
INTERCONNECT DFFT_40_state1_buf_DFFT_44__PIPL_n77(net140_c1,net140);
INTERCONNECT DFFT_41_state2_buf_DFFT_45__PIPL_n78(net141_c1,net141);
INTERCONNECT DFFT_42_state3_buf_DFFT_46__PIPL_n79(net142_c1,net142);
INTERCONNECT SplitCLK_0_211_SplitCLK_0_125(net143_c1,net143);
INTERCONNECT SplitCLK_0_211_SplitCLK_2_166(net144_c1,net144);
INTERCONNECT SplitCLK_4_210_DFFT_78__FPB_n225(net145_c1,net145);
INTERCONNECT SplitCLK_2_209_DFFT_86__FPB_n233(net146_c1,net146);
INTERCONNECT SplitCLK_2_208_DFFT_76__FPB_n223(net147_c1,net147);
INTERCONNECT SplitCLK_2_207_DFFT_84__FPB_n231(net148_c1,net148);
INTERCONNECT SplitCLK_2_206_DFFT_59__FPB_n206(net149_c1,net149);
INTERCONNECT SplitCLK_4_205_DFFT_67__FPB_n214(net150_c1,net150);
INTERCONNECT SplitCLK_4_204_DFFT_75__FPB_n222(net151_c1,net151);
INTERCONNECT SplitCLK_2_203_DFFT_81__FPB_n228(net152_c1,net152);
INTERCONNECT SplitCLK_2_202_DFFT_57__FPB_n204(net153_c1,net153);
INTERCONNECT SplitCLK_4_201_DFFT_65__FPB_n212(net154_c1,net154);
INTERCONNECT SplitCLK_2_200_DFFT_73__FPB_n220(net155_c1,net155);
INTERCONNECT SplitCLK_4_199_DFFT_72__FPB_n219(net156_c1,net156);
INTERCONNECT SplitCLK_2_198_DFFT_80__FPB_n227(net157_c1,net157);
INTERCONNECT SplitCLK_2_197_DFFT_56__FPB_n203(net158_c1,net158);
INTERCONNECT SplitCLK_2_196_DFFT_64__FPB_n211(net159_c1,net159);
INTERCONNECT SplitCLK_2_195_DFFT_55__FPB_n202(net160_c1,net160);
INTERCONNECT SplitCLK_2_194_DFFT_63__FPB_n210(net161_c1,net161);
INTERCONNECT SplitCLK_4_193_DFFT_45__PIPL_n78(net162_c1,net162);
INTERCONNECT SplitCLK_2_192_DFFT_70__FPB_n217(net163_c1,net163);
INTERCONNECT SplitCLK_4_191_DFFT_60__FPB_n207(net164_c1,net164);
INTERCONNECT SplitCLK_4_190_DFFT_51__FBL_n198(net165_c1,net165);
INTERCONNECT SplitCLK_4_189_DFFT_42_state3_buf(net166_c1,net166);
INTERCONNECT SplitCLK_2_188_DFFT_49__ADJFBL_n196(net167_c1,net167);
INTERCONNECT SplitCLK_4_187_DFFT_48__ADJFBL_n195(net168_c1,net168);
INTERCONNECT SplitCLK_4_186_NOTT_16_n40(net169_c1,net169);
INTERCONNECT SplitCLK_4_185_NOTT_14_n38(net170_c1,net170);
INTERCONNECT SplitCLK_4_184_NOTT_10_n34(net171_c1,net171);
INTERCONNECT SplitCLK_4_183_DFFT_40_state1_buf(net172_c1,net172);
INTERCONNECT SplitCLK_4_182_DFFT_47__ADJFBL_n194(net173_c1,net173);
INTERCONNECT SplitCLK_4_181_OR2T_24_n48(net174_c1,net174);
INTERCONNECT SplitCLK_2_180_OR2T_15_n39(net175_c1,net175);
INTERCONNECT SplitCLK_2_179_OR2T_13_n37(net176_c1,net176);
INTERCONNECT SplitCLK_2_178_OR2T_21_n45(net177_c1,net177);
INTERCONNECT SplitCLK_2_177_DFFT_79_state_obs0(net178_c1,net178);
INTERCONNECT SplitCLK_4_176_AND2T_38_n62(net179_c1,net179);
INTERCONNECT SplitCLK_2_175_AND2T_29_n53(net180_c1,net180);
INTERCONNECT SplitCLK_4_174_AND2T_36_n60(net181_c1,net181);
INTERCONNECT SplitCLK_2_173_AND2T_26_n50(net182_c1,net182);
INTERCONNECT SplitCLK_4_172_AND2T_25_n49(net183_c1,net183);
INTERCONNECT SplitCLK_2_171_AND2T_32_n56(net184_c1,net184);
INTERCONNECT SplitCLK_4_170_AND2T_12_n36(net185_c1,net185);
INTERCONNECT SplitCLK_4_169_DFFT_39_state0_buf(net186_c1,net186);
INTERCONNECT SplitCLK_2_168_NOTT_9_n33(net187_c1,net187);
INTERCONNECT SplitCLK_2_167_NOTT_8_n32(net188_c1,net188);
INTERCONNECT SplitCLK_2_166_SplitCLK_6_145(net189_c1,net189);
INTERCONNECT SplitCLK_2_166_SplitCLK_4_165(net190_c1,net190);
INTERCONNECT SplitCLK_4_165_SplitCLK_0_155(net191_c1,net191);
INTERCONNECT SplitCLK_4_165_SplitCLK_2_164(net192_c1,net192);
INTERCONNECT SplitCLK_2_164_SplitCLK_6_159(net193_c1,net193);
INTERCONNECT SplitCLK_2_164_SplitCLK_4_163(net194_c1,net194);
INTERCONNECT SplitCLK_4_163_SplitCLK_2_161(net195_c1,net195);
INTERCONNECT SplitCLK_4_163_SplitCLK_6_162(net196_c1,net196);
INTERCONNECT SplitCLK_6_162_SplitCLK_2_179(net197_c1,net197);
INTERCONNECT SplitCLK_6_162_SplitCLK_4_191(net198_c1,net198);
INTERCONNECT SplitCLK_2_161_SplitCLK_2_206(net199_c1,net199);
INTERCONNECT SplitCLK_2_161_SplitCLK_4_160(net200_c1,net200);
INTERCONNECT SplitCLK_4_160_AND2T_20_n44(net201_c1,net201);
INTERCONNECT SplitCLK_4_160_DFFT_58__FPB_n205(net202_c1,net202);
INTERCONNECT SplitCLK_6_159_SplitCLK_4_157(net203_c1,net203);
INTERCONNECT SplitCLK_6_159_SplitCLK_6_158(net204_c1,net204);
INTERCONNECT SplitCLK_6_158_SplitCLK_2_168(net205_c1,net205);
INTERCONNECT SplitCLK_6_158_SplitCLK_4_201(net206_c1,net206);
INTERCONNECT SplitCLK_4_157_SplitCLK_4_170(net207_c1,net207);
INTERCONNECT SplitCLK_4_157_SplitCLK_4_156(net208_c1,net208);
INTERCONNECT SplitCLK_4_156_AND2T_23_n47(net209_c1,net209);
INTERCONNECT SplitCLK_4_156_OR2T_22_n46(net210_c1,net210);
INTERCONNECT SplitCLK_0_155_SplitCLK_4_150(net211_c1,net211);
INTERCONNECT SplitCLK_0_155_SplitCLK_4_154(net212_c1,net212);
INTERCONNECT SplitCLK_4_154_SplitCLK_0_152(net213_c1,net213);
INTERCONNECT SplitCLK_4_154_SplitCLK_4_153(net214_c1,net214);
INTERCONNECT SplitCLK_4_153_SplitCLK_2_195(net215_c1,net215);
INTERCONNECT SplitCLK_4_153_SplitCLK_2_202(net216_c1,net216);
INTERCONNECT SplitCLK_0_152_SplitCLK_4_176(net217_c1,net217);
INTERCONNECT SplitCLK_0_152_SplitCLK_4_151(net218_c1,net218);
INTERCONNECT SplitCLK_4_151_OR2T_34_n58(net219_c1,net219);
INTERCONNECT SplitCLK_4_151_DFFT_50__FBL_n197(net220_c1,net220);
INTERCONNECT SplitCLK_4_150_SplitCLK_2_147(net221_c1,net221);
INTERCONNECT SplitCLK_4_150_SplitCLK_2_149(net222_c1,net222);
INTERCONNECT SplitCLK_2_149_SplitCLK_2_178(net223_c1,net223);
INTERCONNECT SplitCLK_2_149_SplitCLK_0_148(net224_c1,net224);
INTERCONNECT SplitCLK_0_148_AND2T_27_n51(net225_c1,net225);
INTERCONNECT SplitCLK_0_148_DFFT_61__FPB_n208(net226_c1,net226);
INTERCONNECT SplitCLK_2_147_SplitCLK_2_180(net227_c1,net227);
INTERCONNECT SplitCLK_2_147_SplitCLK_4_146(net228_c1,net228);
INTERCONNECT SplitCLK_4_146_XOR2T_28_n52(net229_c1,net229);
INTERCONNECT SplitCLK_4_146_OR2T_11_n35(net230_c1,net230);
INTERCONNECT SplitCLK_6_145_SplitCLK_4_135(net231_c1,net231);
INTERCONNECT SplitCLK_6_145_SplitCLK_6_144(net232_c1,net232);
INTERCONNECT SplitCLK_6_144_SplitCLK_6_139(net233_c1,net233);
INTERCONNECT SplitCLK_6_144_SplitCLK_4_143(net234_c1,net234);
INTERCONNECT SplitCLK_4_143_SplitCLK_4_141(net235_c1,net235);
INTERCONNECT SplitCLK_4_143_SplitCLK_6_142(net236_c1,net236);
INTERCONNECT SplitCLK_6_142_SplitCLK_4_182(net237_c1,net237);
INTERCONNECT SplitCLK_6_142_SplitCLK_2_208(net238_c1,net238);
INTERCONNECT SplitCLK_4_141_SplitCLK_4_190(net239_c1,net239);
INTERCONNECT SplitCLK_4_141_SplitCLK_4_140(net240_c1,net240);
INTERCONNECT SplitCLK_4_140_DFFT_52__FBL_n199(net241_c1,net241);
INTERCONNECT SplitCLK_4_140_DFFT_43__PIPL_n76(net242_c1,net242);
INTERCONNECT SplitCLK_6_139_SplitCLK_0_137(net243_c1,net243);
INTERCONNECT SplitCLK_6_139_SplitCLK_6_138(net244_c1,net244);
INTERCONNECT SplitCLK_6_138_SplitCLK_2_177(net245_c1,net245);
INTERCONNECT SplitCLK_6_138_SplitCLK_4_210(net246_c1,net246);
INTERCONNECT SplitCLK_0_137_SplitCLK_4_169(net247_c1,net247);
INTERCONNECT SplitCLK_0_137_SplitCLK_4_136(net248_c1,net248);
INTERCONNECT SplitCLK_4_136_DFFT_83_state_obs1(net249_c1,net249);
INTERCONNECT SplitCLK_4_136_DFFT_77__FPB_n224(net250_c1,net250);
INTERCONNECT SplitCLK_4_135_SplitCLK_6_130(net251_c1,net251);
INTERCONNECT SplitCLK_4_135_SplitCLK_0_134(net252_c1,net252);
INTERCONNECT SplitCLK_0_134_SplitCLK_4_132(net253_c1,net253);
INTERCONNECT SplitCLK_0_134_SplitCLK_2_133(net254_c1,net254);
INTERCONNECT SplitCLK_2_133_SplitCLK_4_187(net255_c1,net255);
INTERCONNECT SplitCLK_2_133_SplitCLK_2_203(net256_c1,net256);
INTERCONNECT SplitCLK_4_132_SplitCLK_2_175(net257_c1,net257);
INTERCONNECT SplitCLK_4_132_SplitCLK_4_131(net258_c1,net258);
INTERCONNECT SplitCLK_4_131_OR2T_30_n54(net259_c1,net259);
INTERCONNECT SplitCLK_4_131_DFFT_66__FPB_n213(net260_c1,net260);
INTERCONNECT SplitCLK_6_130_SplitCLK_0_127(net261_c1,net261);
INTERCONNECT SplitCLK_6_130_SplitCLK_2_129(net262_c1,net262);
INTERCONNECT SplitCLK_2_129_SplitCLK_2_198(net263_c1,net263);
INTERCONNECT SplitCLK_2_129_SplitCLK_4_128(net264_c1,net264);
INTERCONNECT SplitCLK_4_128_DFFT_44__PIPL_n77(net265_c1,net265);
INTERCONNECT SplitCLK_4_128_DFFT_82__FPB_n229(net266_c1,net266);
INTERCONNECT SplitCLK_0_127_SplitCLK_4_183(net267_c1,net267);
INTERCONNECT SplitCLK_0_127_SplitCLK_0_126(net268_c1,net268);
INTERCONNECT SplitCLK_0_126_DFFT_87_state_obs2(net269_c1,net269);
INTERCONNECT SplitCLK_0_126_DFFT_85__FPB_n232(net270_c1,net270);
INTERCONNECT SplitCLK_0_125_SplitCLK_6_104(net271_c1,net271);
INTERCONNECT SplitCLK_0_125_SplitCLK_4_124(net272_c1,net272);
INTERCONNECT SplitCLK_4_124_SplitCLK_0_114(net273_c1,net273);
INTERCONNECT SplitCLK_4_124_SplitCLK_2_123(net274_c1,net274);
INTERCONNECT SplitCLK_2_123_SplitCLK_6_118(net275_c1,net275);
INTERCONNECT SplitCLK_2_123_SplitCLK_4_122(net276_c1,net276);
INTERCONNECT SplitCLK_4_122_SplitCLK_4_120(net277_c1,net277);
INTERCONNECT SplitCLK_4_122_SplitCLK_2_121(net278_c1,net278);
INTERCONNECT SplitCLK_2_121_SplitCLK_2_200(net279_c1,net279);
INTERCONNECT SplitCLK_2_121_SplitCLK_4_204(net280_c1,net280);
INTERCONNECT SplitCLK_4_120_SplitCLK_4_174(net281_c1,net281);
INTERCONNECT SplitCLK_4_120_SplitCLK_4_119(net282_c1,net282);
INTERCONNECT SplitCLK_4_119_AND2T_19_n43(net283_c1,net283);
INTERCONNECT SplitCLK_4_119_AND2T_37_n61(net284_c1,net284);
INTERCONNECT SplitCLK_6_118_SplitCLK_0_116(net285_c1,net285);
INTERCONNECT SplitCLK_6_118_SplitCLK_6_117(net286_c1,net286);
INTERCONNECT SplitCLK_6_117_SplitCLK_4_172(net287_c1,net287);
INTERCONNECT SplitCLK_6_117_SplitCLK_2_173(net288_c1,net288);
INTERCONNECT SplitCLK_0_116_SplitCLK_4_181(net289_c1,net289);
INTERCONNECT SplitCLK_0_116_SplitCLK_4_115(net290_c1,net290);
INTERCONNECT SplitCLK_4_115_OR2T_35_n59(net291_c1,net291);
INTERCONNECT SplitCLK_4_115_DFFT_74__FPB_n221(net292_c1,net292);
INTERCONNECT SplitCLK_0_114_SplitCLK_4_109(net293_c1,net293);
INTERCONNECT SplitCLK_0_114_SplitCLK_4_113(net294_c1,net294);
INTERCONNECT SplitCLK_4_113_SplitCLK_0_111(net295_c1,net295);
INTERCONNECT SplitCLK_4_113_SplitCLK_4_112(net296_c1,net296);
INTERCONNECT SplitCLK_4_112_SplitCLK_2_194(net297_c1,net297);
INTERCONNECT SplitCLK_4_112_SplitCLK_2_196(net298_c1,net298);
INTERCONNECT SplitCLK_0_111_SplitCLK_4_185(net299_c1,net299);
INTERCONNECT SplitCLK_0_111_SplitCLK_4_110(net300_c1,net300);
INTERCONNECT SplitCLK_4_110_DFFT_71__FPB_n218(net301_c1,net301);
INTERCONNECT SplitCLK_4_110_DFFT_68__FPB_n215(net302_c1,net302);
INTERCONNECT SplitCLK_4_109_SplitCLK_4_106(net303_c1,net303);
INTERCONNECT SplitCLK_4_109_SplitCLK_2_108(net304_c1,net304);
INTERCONNECT SplitCLK_2_108_SplitCLK_2_167(net305_c1,net305);
INTERCONNECT SplitCLK_2_108_SplitCLK_4_107(net306_c1,net306);
INTERCONNECT SplitCLK_4_107_OR2T_18_n42(net307_c1,net307);
INTERCONNECT SplitCLK_4_107_DFFT_62__FPB_n209(net308_c1,net308);
INTERCONNECT SplitCLK_4_106_SplitCLK_4_205(net309_c1,net309);
INTERCONNECT SplitCLK_4_106_SplitCLK_4_105(net310_c1,net310);
INTERCONNECT SplitCLK_4_105_OR2T_17_n41(net311_c1,net311);
INTERCONNECT SplitCLK_4_105_DFFT_69__FPB_n216(net312_c1,net312);
INTERCONNECT SplitCLK_6_104_SplitCLK_6_94(net313_c1,net313);
INTERCONNECT SplitCLK_6_104_SplitCLK_6_103(net314_c1,net314);
INTERCONNECT SplitCLK_6_103_SplitCLK_6_98(net315_c1,net315);
INTERCONNECT SplitCLK_6_103_SplitCLK_4_102(net316_c1,net316);
INTERCONNECT SplitCLK_4_102_SplitCLK_4_100(net317_c1,net317);
INTERCONNECT SplitCLK_4_102_SplitCLK_6_101(net318_c1,net318);
INTERCONNECT SplitCLK_6_101_SplitCLK_2_192(net319_c1,net319);
INTERCONNECT SplitCLK_6_101_SplitCLK_4_199(net320_c1,net320);
INTERCONNECT SplitCLK_4_100_SplitCLK_4_184(net321_c1,net321);
INTERCONNECT SplitCLK_4_100_SplitCLK_4_99(net322_c1,net322);
INTERCONNECT SplitCLK_4_99_OR2T_31_n55(net323_c1,net323);
INTERCONNECT SplitCLK_4_99_DFFT_53__FBL_n200(net324_c1,net324);
INTERCONNECT SplitCLK_6_98_SplitCLK_2_96(net325_c1,net325);
INTERCONNECT SplitCLK_6_98_SplitCLK_6_97(net326_c1,net326);
INTERCONNECT SplitCLK_6_97_SplitCLK_4_193(net327_c1,net327);
INTERCONNECT SplitCLK_6_97_SplitCLK_2_209(net328_c1,net328);
INTERCONNECT SplitCLK_2_96_SplitCLK_2_207(net329_c1,net329);
INTERCONNECT SplitCLK_2_96_SplitCLK_4_95(net330_c1,net330);
INTERCONNECT SplitCLK_4_95_DFFT_91_state_obs3(net331_c1,net331);
INTERCONNECT SplitCLK_4_95_DFFT_41_state2_buf(net332_c1,net332);
INTERCONNECT SplitCLK_6_94_SplitCLK_4_89(net333_c1,net333);
INTERCONNECT SplitCLK_6_94_SplitCLK_4_93(net334_c1,net334);
INTERCONNECT SplitCLK_4_93_SplitCLK_0_91(net335_c1,net335);
INTERCONNECT SplitCLK_4_93_SplitCLK_4_92(net336_c1,net336);
INTERCONNECT SplitCLK_4_92_SplitCLK_2_171(net337_c1,net337);
INTERCONNECT SplitCLK_4_92_SplitCLK_2_197(net338_c1,net338);
INTERCONNECT SplitCLK_0_91_SplitCLK_4_186(net339_c1,net339);
INTERCONNECT SplitCLK_0_91_SplitCLK_4_90(net340_c1,net340);
INTERCONNECT SplitCLK_4_90_AND2T_33_n57(net341_c1,net341);
INTERCONNECT SplitCLK_4_90_DFFT_54__FPB_n201(net342_c1,net342);
INTERCONNECT SplitCLK_4_89_SplitCLK_4_86(net343_c1,net343);
INTERCONNECT SplitCLK_4_89_SplitCLK_6_88(net344_c1,net344);
INTERCONNECT SplitCLK_6_88_SplitCLK_2_188(net345_c1,net345);
INTERCONNECT SplitCLK_6_88_SplitCLK_4_87(net346_c1,net346);
INTERCONNECT SplitCLK_4_87_DFFT_46__PIPL_n79(net347_c1,net347);
INTERCONNECT SplitCLK_4_87_DFFT_88__FPB_n235(net348_c1,net348);
INTERCONNECT SplitCLK_4_86_SplitCLK_4_189(net349_c1,net349);
INTERCONNECT SplitCLK_4_86_SplitCLK_4_85(net350_c1,net350);
INTERCONNECT SplitCLK_4_85_DFFT_90__FPB_n237(net351_c1,net351);
INTERCONNECT SplitCLK_4_85_DFFT_89__FPB_n236(net352_c1,net352);
INTERCONNECT GCLK_Pad_SplitCLK_0_211(GCLK_Pad,net353);

endmodule
