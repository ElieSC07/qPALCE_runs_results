module KSA4_route(
input GCLK_Pad,
input a0_Pad,
input a1_Pad,
input b0_Pad,
input a2_Pad,
input b1_Pad,
input a3_Pad,
input b2_Pad,
input b3_Pad,
input cin_Pad,
output cout_Pad,
output sum0_Pad,
output sum1_Pad,
output sum2_Pad,
output sum3_Pad);

wire a0_Pad;
wire net0;
wire a1_Pad;
wire net1;
wire b0_Pad;
wire net2;
wire a2_Pad;
wire net3;
wire b1_Pad;
wire net4;
wire a3_Pad;
wire net5;
wire b2_Pad;
wire net6;
wire b3_Pad;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire cin_Pad;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire cout_Pad;
wire net66_c1;
wire sum0_Pad;
wire net67_c1;
wire sum1_Pad;
wire net68_c1;
wire sum2_Pad;
wire net69_c1;
wire sum3_Pad;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire GCLK_Pad;
wire net247;

XOR2T XOR2T_21_n21(net155,net79,net97,net9_c1);
XOR2T XOR2T_30_n30(net245,net74,net88,net10_c1);
XOR2T XOR2T_22_n22(net229,net72,net85,net11_c1);
XOR2T XOR2T_15_n15(net169,net70,net77,net14_c1);
XOR2T XOR2T_16_n16(net149,net89,net106,net18_c1);
XOR2T XOR2T_17_n17(net185,net71,net81,net22_c1);
XOR2T XOR2T_29_n29(net215,net33,net112,net34_c1);
XOR2T XOR2T_37_sum3(net239,net32,net109,net69_c1);
AND2T AND2T_31_n31(net223,net87,net73,net12_c1);
AND2T AND2T_23_n23(net151,net93,net86,net13_c1);
AND2T AND2T_40_n40(net207,net60,net116,net15_c1);
AND2T AND2T_32_n32(net225,net46,net117,net16_c1);
AND2T AND2T_24_n24(net157,net13,net100,net17_c1);
AND2T AND2T_41_n41(net177,net80,net45,net19_c1);
AND2T AND2T_33_n33(net171,net94,net53,net20_c1);
AND2T AND2T_25_n25(net165,net75,net62,net21_c1);
AND2T AND2T_42_n42(net230,net42,net57,net23_c1);
AND2T AND2T_34_n34(net231,net41,net55,net24_c1);
AND2T AND2T_26_n26(net183,net39,net51,net25_c1);
AND2T AND2T_18_n18(net143,net58,net110,net26_c1);
AND2T AND2T_19_n19(net170,net38,net47,net30_c1);
AND2T AND2T_38_n38(net232,net76,net90,net35_c1);
AND2T AND2T_39_n39(net199,net63,net111,net36_c1);
OR2T OR2T_20_n20(net144,net26,net113,net8_c1);
OR2T OR2T_43_n43(net184,net19,net118,net27_c1);
OR2T OR2T_35_n35(net178,net20,net119,net28_c1);
OR2T OR2T_27_n27(net166,net21,net102,net29_c1);
OR2T OR2T_44_n44(net158,net15,net120,net31_c1);
OR2T OR2T_36_n36(net240,net16,net121,net32_c1);
OR2T OR2T_28_n28(net209,net95,net92,net33_c1);
DFFT DFFT_72_sum0(net128,net107,net66_c1);
DFFT DFFT_74_sum1(net195,net114,net67_c1);
DFFT DFFT_75_sum2(net210,net34,net68_c1);
DFFT DFFT_50__FPB_n140(net156,net115,net97_c1);
DFFT DFFT_51__FPB_n141(net137,net78,net98_c1);
DFFT DFFT_60__FPB_n150(net243,net96,net99_c1);
DFFT DFFT_52__FPB_n142(net127,net98,net100_c1);
OR2T OR2T_45_cout(net200,net31,net122,net65_c1);
DFFT DFFT_61__FPB_n151(net237,net99,net101_c1);
DFFT DFFT_53__FPB_n143(net126,net61,net102_c1);
DFFT DFFT_70__FPB_n160(net152,net123,net103_c1);
DFFT DFFT_62__FPB_n152(net244,net101,net104_c1);
DFFT DFFT_54__FPB_n144(net238,net56,net105_c1);
DFFT DFFT_46__FPB_n136(net138,net82,net106_c1);
DFFT DFFT_71__FPB_n161(net196,net103,net107_c1);
DFFT DFFT_63__FPB_n153(net246,net104,net109_c1);
DFFT DFFT_55__FPB_n145(net213,net105,net108_c1);
DFFT DFFT_47__FPB_n137(net141,net49,net110_c1);
DFFT DFFT_64__FPB_n154(net201,net84,net111_c1);
DFFT DFFT_56__FPB_n146(net214,net108,net112_c1);
DFFT DFFT_48__FPB_n138(net142,net43,net113_c1);
DFFT DFFT_73__FPB_n163(net208,net9,net114_c1);
DFFT DFFT_65__FPB_n155(net216,net52,net116_c1);
DFFT DFFT_57__FPB_n147(net226,net12,net117_c1);
DFFT DFFT_49__FPB_n139(net179,net40,net115_c1);
DFFT DFFT_66__FPB_n156(net186,net23,net118_c1);
DFFT DFFT_58__FPB_n148(net172,net50,net119_c1);
SPLITT Split_100_n190(net64,net45_c1,net76_c1);
SPLITT Split_101_n191(net24,net50_c1,net80_c1);
SPLITT Split_102_n192(net35,net52_c1,net84_c1);
DFFT DFFT_67__FPB_n157(net224,net27,net120_c1);
DFFT DFFT_59__FPB_n149(net180,net28,net121_c1);
DFFT DFFT_68__FPB_n158(net202,net36,net122_c1);
DFFT DFFT_69__FPB_n159(net150,net18,net123_c1);
SPLITT Split_80_n170(net2,net38_c1,net70_c1);
SPLITT Split_81_n171(net4,net39_c1,net71_c1);
SPLITT Split_82_n172(net6,net41_c1,net72_c1);
SPLITT Split_90_n180(net59,net40_c1,net73_c1);
SPLITT Split_83_n173(net7,net42_c1,net74_c1);
SPLITT Split_91_n181(net30,net43_c1,net75_c1);
SPLITT Split_76_n166(net0,net47_c1,net77_c1);
SPLITT Split_84_n174(net37,net44_c1,net78_c1);
SPLITT Split_92_n182(net8,net46_c1,net79_c1);
SPLITT Split_77_n167(net1,net51_c1,net81_c1);
SPLITT Split_85_n175(net44,net49_c1,net82_c1);
SPLITT Split_93_n183(net11,net48_c1,net83_c1);
SPLITT Split_78_n168(net3,net55_c1,net85_c1);
SPLITT Split_86_n176(net14,net54_c1,net86_c1);
SPLITT Split_94_n184(net83,net53_c1,net87_c1);
SPLITT Split_79_n169(net5,net57_c1,net88_c1);
SPLITT Split_87_n177(net54,net58_c1,net89_c1);
SPLITT Split_95_n185(net48,net56_c1,net90_c1);
SPLITT Split_88_n178(net22,net59_c1,net91_c1);
SPLITT Split_96_n186(net17,net60_c1,net92_c1);
SPLITT Split_89_n179(net91,net62_c1,net93_c1);
SPLITT Split_97_n187(net25,net61_c1,net94_c1);
SPLITT Split_98_n188(net29,net63_c1,net95_c1);
SPLITT Split_99_n189(net10,net64_c1,net96_c1);
SPLITT SplitCLK_4_62(net241,net245_c1,net246_c1);
SPLITT SplitCLK_4_63(net242,net243_c1,net244_c1);
SPLITT SplitCLK_6_64(net233,net241_c1,net242_c1);
SPLITT SplitCLK_4_65(net235,net240_c1,net239_c1);
SPLITT SplitCLK_4_66(net236,net237_c1,net238_c1);
SPLITT SplitCLK_4_67(net234,net236_c1,net235_c1);
SPLITT SplitCLK_0_68(net217,net233_c1,net234_c1);
SPLITT SplitCLK_4_69(net227,net232_c1,net231_c1);
SPLITT SplitCLK_4_70(net228,net230_c1,net229_c1);
SPLITT SplitCLK_6_71(net219,net227_c1,net228_c1);
SPLITT SplitCLK_4_72(net221,net226_c1,net225_c1);
SPLITT SplitCLK_4_73(net222,net224_c1,net223_c1);
SPLITT SplitCLK_2_74(net220,net221_c1,net222_c1);
SPLITT SplitCLK_6_75(net218,net219_c1,net220_c1);
SPLITT SplitCLK_2_76(net187,net217_c1,net218_c1);
SPLITT SplitCLK_4_77(net211,net215_c1,net216_c1);
SPLITT SplitCLK_4_78(net212,net213_c1,net214_c1);
SPLITT SplitCLK_4_79(net203,net212_c1,net211_c1);
SPLITT SplitCLK_4_80(net205,net209_c1,net210_c1);
SPLITT SplitCLK_4_81(net206,net207_c1,net208_c1);
SPLITT SplitCLK_4_82(net204,net206_c1,net205_c1);
SPLITT SplitCLK_0_83(net189,net203_c1,net204_c1);
SPLITT SplitCLK_4_84(net197,net201_c1,net202_c1);
SPLITT SplitCLK_4_85(net198,net199_c1,net200_c1);
SPLITT SplitCLK_6_86(net191,net197_c1,net198_c1);
SPLITT SplitCLK_4_87(net194,net196_c1,net195_c1);
SPLITT SplitCLK_4_88(net192,net193_c1,net194_c1);
SPLITT SplitCLK_4_89(net190,net191_c1,net192_c1);
SPLITT SplitCLK_4_90(net188,net190_c1,net189_c1);
SPLITT SplitCLK_0_91(net124,net187_c1,net188_c1);
SPLITT SplitCLK_4_92(net181,net185_c1,net186_c1);
SPLITT SplitCLK_4_93(net182,net183_c1,net184_c1);
SPLITT SplitCLK_4_94(net173,net182_c1,net181_c1);
SPLITT SplitCLK_4_95(net175,net180_c1,net179_c1);
SPLITT SplitCLK_4_96(net176,net177_c1,net178_c1);
SPLITT SplitCLK_4_97(net174,net176_c1,net175_c1);
SPLITT SplitCLK_4_98(net159,net173_c1,net174_c1);
SPLITT SplitCLK_4_99(net167,net172_c1,net171_c1);
SPLITT SplitCLK_4_100(net168,net170_c1,net169_c1);
SPLITT SplitCLK_2_101(net161,net167_c1,net168_c1);
SPLITT SplitCLK_4_102(net164,net165_c1,net166_c1);
SPLITT SplitCLK_4_103(net162,net163_c1,net164_c1);
SPLITT SplitCLK_2_104(net160,net162_c1,net161_c1);
SPLITT SplitCLK_6_105(net129,net159_c1,net160_c1);
SPLITT SplitCLK_4_106(net153,net158_c1,net157_c1);
SPLITT SplitCLK_0_107(net154,net155_c1,net156_c1);
SPLITT SplitCLK_6_108(net145,net153_c1,net154_c1);
SPLITT SplitCLK_4_109(net147,net151_c1,net152_c1);
SPLITT SplitCLK_4_110(net148,net149_c1,net150_c1);
SPLITT SplitCLK_4_111(net146,net148_c1,net147_c1);
SPLITT SplitCLK_4_112(net131,net145_c1,net146_c1);
SPLITT SplitCLK_4_113(net139,net144_c1,net143_c1);
SPLITT SplitCLK_4_114(net140,net142_c1,net141_c1);
SPLITT SplitCLK_2_115(net133,net139_c1,net140_c1);
SPLITT SplitCLK_4_116(net136,net137_c1,net138_c1);
SPLITT SplitCLK_4_117(net134,net135_c1,net136_c1);
SPLITT SplitCLK_6_118(net132,net134_c1,net133_c1);
SPLITT SplitCLK_4_119(net130,net132_c1,net131_c1);
SPLITT SplitCLK_2_120(net125,net130_c1,net129_c1);
wire dummy0;
SPLITT SplitCLK_2_121(net193,net128_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_2_122(net135,net127_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_123(net163,net126_c1,dummy2);
SPLITT SplitCLK_0_124(net247,net124_c1,net125_c1);
INTERCONNECT a0_Pad_Split_76_n166(a0_Pad,net0);
INTERCONNECT a1_Pad_Split_77_n167(a1_Pad,net1);
INTERCONNECT b0_Pad_Split_80_n170(b0_Pad,net2);
INTERCONNECT a2_Pad_Split_78_n168(a2_Pad,net3);
INTERCONNECT b1_Pad_Split_81_n171(b1_Pad,net4);
INTERCONNECT a3_Pad_Split_79_n169(a3_Pad,net5);
INTERCONNECT b2_Pad_Split_82_n172(b2_Pad,net6);
INTERCONNECT b3_Pad_Split_83_n173(b3_Pad,net7);
INTERCONNECT OR2T_20_n20_Split_92_n182(net8_c1,net8);
INTERCONNECT XOR2T_21_n21_DFFT_73__FPB_n163(net9_c1,net9);
INTERCONNECT XOR2T_30_n30_Split_99_n189(net10_c1,net10);
INTERCONNECT XOR2T_22_n22_Split_93_n183(net11_c1,net11);
INTERCONNECT AND2T_31_n31_DFFT_57__FPB_n147(net12_c1,net12);
INTERCONNECT AND2T_23_n23_AND2T_24_n24(net13_c1,net13);
INTERCONNECT XOR2T_15_n15_Split_86_n176(net14_c1,net14);
INTERCONNECT AND2T_40_n40_OR2T_44_n44(net15_c1,net15);
INTERCONNECT AND2T_32_n32_OR2T_36_n36(net16_c1,net16);
INTERCONNECT AND2T_24_n24_Split_96_n186(net17_c1,net17);
INTERCONNECT XOR2T_16_n16_DFFT_69__FPB_n159(net18_c1,net18);
INTERCONNECT AND2T_41_n41_OR2T_43_n43(net19_c1,net19);
INTERCONNECT AND2T_33_n33_OR2T_35_n35(net20_c1,net20);
INTERCONNECT AND2T_25_n25_OR2T_27_n27(net21_c1,net21);
INTERCONNECT XOR2T_17_n17_Split_88_n178(net22_c1,net22);
INTERCONNECT AND2T_42_n42_DFFT_66__FPB_n156(net23_c1,net23);
INTERCONNECT AND2T_34_n34_Split_101_n191(net24_c1,net24);
INTERCONNECT AND2T_26_n26_Split_97_n187(net25_c1,net25);
INTERCONNECT AND2T_18_n18_OR2T_20_n20(net26_c1,net26);
INTERCONNECT OR2T_43_n43_DFFT_67__FPB_n157(net27_c1,net27);
INTERCONNECT OR2T_35_n35_DFFT_59__FPB_n149(net28_c1,net28);
INTERCONNECT OR2T_27_n27_Split_98_n188(net29_c1,net29);
INTERCONNECT AND2T_19_n19_Split_91_n181(net30_c1,net30);
INTERCONNECT OR2T_44_n44_OR2T_45_cout(net31_c1,net31);
INTERCONNECT OR2T_36_n36_XOR2T_37_sum3(net32_c1,net32);
INTERCONNECT OR2T_28_n28_XOR2T_29_n29(net33_c1,net33);
INTERCONNECT XOR2T_29_n29_DFFT_75_sum2(net34_c1,net34);
INTERCONNECT AND2T_38_n38_Split_102_n192(net35_c1,net35);
INTERCONNECT AND2T_39_n39_DFFT_68__FPB_n158(net36_c1,net36);
INTERCONNECT cin_Pad_Split_84_n174(cin_Pad,net37);
INTERCONNECT Split_80_n170_AND2T_19_n19(net38_c1,net38);
INTERCONNECT Split_81_n171_AND2T_26_n26(net39_c1,net39);
INTERCONNECT Split_90_n180_DFFT_49__FPB_n139(net40_c1,net40);
INTERCONNECT Split_82_n172_AND2T_34_n34(net41_c1,net41);
INTERCONNECT Split_83_n173_AND2T_42_n42(net42_c1,net42);
INTERCONNECT Split_91_n181_DFFT_48__FPB_n138(net43_c1,net43);
INTERCONNECT Split_84_n174_Split_85_n175(net44_c1,net44);
INTERCONNECT Split_100_n190_AND2T_41_n41(net45_c1,net45);
INTERCONNECT Split_92_n182_AND2T_32_n32(net46_c1,net46);
INTERCONNECT Split_76_n166_AND2T_19_n19(net47_c1,net47);
INTERCONNECT Split_93_n183_Split_95_n185(net48_c1,net48);
INTERCONNECT Split_85_n175_DFFT_47__FPB_n137(net49_c1,net49);
INTERCONNECT Split_101_n191_DFFT_58__FPB_n148(net50_c1,net50);
INTERCONNECT Split_77_n167_AND2T_26_n26(net51_c1,net51);
INTERCONNECT Split_102_n192_DFFT_65__FPB_n155(net52_c1,net52);
INTERCONNECT Split_94_n184_AND2T_33_n33(net53_c1,net53);
INTERCONNECT Split_86_n176_Split_87_n177(net54_c1,net54);
INTERCONNECT Split_78_n168_AND2T_34_n34(net55_c1,net55);
INTERCONNECT Split_95_n185_DFFT_54__FPB_n144(net56_c1,net56);
INTERCONNECT Split_79_n169_AND2T_42_n42(net57_c1,net57);
INTERCONNECT Split_87_n177_AND2T_18_n18(net58_c1,net58);
INTERCONNECT Split_88_n178_Split_90_n180(net59_c1,net59);
INTERCONNECT Split_96_n186_AND2T_40_n40(net60_c1,net60);
INTERCONNECT Split_97_n187_DFFT_53__FPB_n143(net61_c1,net61);
INTERCONNECT Split_89_n179_AND2T_25_n25(net62_c1,net62);
INTERCONNECT Split_98_n188_AND2T_39_n39(net63_c1,net63);
INTERCONNECT Split_99_n189_Split_100_n190(net64_c1,net64);
INTERCONNECT OR2T_45_cout_cout_Pad(net65_c1,cout_Pad);
INTERCONNECT DFFT_72_sum0_sum0_Pad(net66_c1,sum0_Pad);
INTERCONNECT DFFT_74_sum1_sum1_Pad(net67_c1,sum1_Pad);
INTERCONNECT DFFT_75_sum2_sum2_Pad(net68_c1,sum2_Pad);
INTERCONNECT XOR2T_37_sum3_sum3_Pad(net69_c1,sum3_Pad);
INTERCONNECT Split_80_n170_XOR2T_15_n15(net70_c1,net70);
INTERCONNECT Split_81_n171_XOR2T_17_n17(net71_c1,net71);
INTERCONNECT Split_82_n172_XOR2T_22_n22(net72_c1,net72);
INTERCONNECT Split_90_n180_AND2T_31_n31(net73_c1,net73);
INTERCONNECT Split_83_n173_XOR2T_30_n30(net74_c1,net74);
INTERCONNECT Split_91_n181_AND2T_25_n25(net75_c1,net75);
INTERCONNECT Split_100_n190_AND2T_38_n38(net76_c1,net76);
INTERCONNECT Split_76_n166_XOR2T_15_n15(net77_c1,net77);
INTERCONNECT Split_84_n174_DFFT_51__FPB_n141(net78_c1,net78);
INTERCONNECT Split_92_n182_XOR2T_21_n21(net79_c1,net79);
INTERCONNECT Split_101_n191_AND2T_41_n41(net80_c1,net80);
INTERCONNECT Split_77_n167_XOR2T_17_n17(net81_c1,net81);
INTERCONNECT Split_85_n175_DFFT_46__FPB_n136(net82_c1,net82);
INTERCONNECT Split_93_n183_Split_94_n184(net83_c1,net83);
INTERCONNECT Split_102_n192_DFFT_64__FPB_n154(net84_c1,net84);
INTERCONNECT Split_78_n168_XOR2T_22_n22(net85_c1,net85);
INTERCONNECT Split_86_n176_AND2T_23_n23(net86_c1,net86);
INTERCONNECT Split_94_n184_AND2T_31_n31(net87_c1,net87);
INTERCONNECT Split_79_n169_XOR2T_30_n30(net88_c1,net88);
INTERCONNECT Split_87_n177_XOR2T_16_n16(net89_c1,net89);
INTERCONNECT Split_95_n185_AND2T_38_n38(net90_c1,net90);
INTERCONNECT Split_88_n178_Split_89_n179(net91_c1,net91);
INTERCONNECT Split_96_n186_OR2T_28_n28(net92_c1,net92);
INTERCONNECT Split_89_n179_AND2T_23_n23(net93_c1,net93);
INTERCONNECT Split_97_n187_AND2T_33_n33(net94_c1,net94);
INTERCONNECT Split_98_n188_OR2T_28_n28(net95_c1,net95);
INTERCONNECT Split_99_n189_DFFT_60__FPB_n150(net96_c1,net96);
INTERCONNECT DFFT_50__FPB_n140_XOR2T_21_n21(net97_c1,net97);
INTERCONNECT DFFT_51__FPB_n141_DFFT_52__FPB_n142(net98_c1,net98);
INTERCONNECT DFFT_60__FPB_n150_DFFT_61__FPB_n151(net99_c1,net99);
INTERCONNECT DFFT_52__FPB_n142_AND2T_24_n24(net100_c1,net100);
INTERCONNECT DFFT_61__FPB_n151_DFFT_62__FPB_n152(net101_c1,net101);
INTERCONNECT DFFT_53__FPB_n143_OR2T_27_n27(net102_c1,net102);
INTERCONNECT DFFT_70__FPB_n160_DFFT_71__FPB_n161(net103_c1,net103);
INTERCONNECT DFFT_62__FPB_n152_DFFT_63__FPB_n153(net104_c1,net104);
INTERCONNECT DFFT_54__FPB_n144_DFFT_55__FPB_n145(net105_c1,net105);
INTERCONNECT DFFT_46__FPB_n136_XOR2T_16_n16(net106_c1,net106);
INTERCONNECT DFFT_71__FPB_n161_DFFT_72_sum0(net107_c1,net107);
INTERCONNECT DFFT_55__FPB_n145_DFFT_56__FPB_n146(net108_c1,net108);
INTERCONNECT DFFT_63__FPB_n153_XOR2T_37_sum3(net109_c1,net109);
INTERCONNECT DFFT_47__FPB_n137_AND2T_18_n18(net110_c1,net110);
INTERCONNECT DFFT_64__FPB_n154_AND2T_39_n39(net111_c1,net111);
INTERCONNECT DFFT_56__FPB_n146_XOR2T_29_n29(net112_c1,net112);
INTERCONNECT DFFT_48__FPB_n138_OR2T_20_n20(net113_c1,net113);
INTERCONNECT DFFT_73__FPB_n163_DFFT_74_sum1(net114_c1,net114);
INTERCONNECT DFFT_49__FPB_n139_DFFT_50__FPB_n140(net115_c1,net115);
INTERCONNECT DFFT_65__FPB_n155_AND2T_40_n40(net116_c1,net116);
INTERCONNECT DFFT_57__FPB_n147_AND2T_32_n32(net117_c1,net117);
INTERCONNECT DFFT_66__FPB_n156_OR2T_43_n43(net118_c1,net118);
INTERCONNECT DFFT_58__FPB_n148_OR2T_35_n35(net119_c1,net119);
INTERCONNECT DFFT_67__FPB_n157_OR2T_44_n44(net120_c1,net120);
INTERCONNECT DFFT_59__FPB_n149_OR2T_36_n36(net121_c1,net121);
INTERCONNECT DFFT_68__FPB_n158_OR2T_45_cout(net122_c1,net122);
INTERCONNECT DFFT_69__FPB_n159_DFFT_70__FPB_n160(net123_c1,net123);
INTERCONNECT SplitCLK_0_124_SplitCLK_0_91(net124_c1,net124);
INTERCONNECT SplitCLK_0_124_SplitCLK_2_120(net125_c1,net125);
INTERCONNECT SplitCLK_2_123_DFFT_53__FPB_n143(net126_c1,net126);
INTERCONNECT SplitCLK_2_122_DFFT_52__FPB_n142(net127_c1,net127);
INTERCONNECT SplitCLK_2_121_DFFT_72_sum0(net128_c1,net128);
INTERCONNECT SplitCLK_2_120_SplitCLK_6_105(net129_c1,net129);
INTERCONNECT SplitCLK_2_120_SplitCLK_4_119(net130_c1,net130);
INTERCONNECT SplitCLK_4_119_SplitCLK_4_112(net131_c1,net131);
INTERCONNECT SplitCLK_4_119_SplitCLK_6_118(net132_c1,net132);
INTERCONNECT SplitCLK_6_118_SplitCLK_2_115(net133_c1,net133);
INTERCONNECT SplitCLK_6_118_SplitCLK_4_117(net134_c1,net134);
INTERCONNECT SplitCLK_4_117_SplitCLK_2_122(net135_c1,net135);
INTERCONNECT SplitCLK_4_117_SplitCLK_4_116(net136_c1,net136);
INTERCONNECT SplitCLK_4_116_DFFT_51__FPB_n141(net137_c1,net137);
INTERCONNECT SplitCLK_4_116_DFFT_46__FPB_n136(net138_c1,net138);
INTERCONNECT SplitCLK_2_115_SplitCLK_4_113(net139_c1,net139);
INTERCONNECT SplitCLK_2_115_SplitCLK_4_114(net140_c1,net140);
INTERCONNECT SplitCLK_4_114_DFFT_47__FPB_n137(net141_c1,net141);
INTERCONNECT SplitCLK_4_114_DFFT_48__FPB_n138(net142_c1,net142);
INTERCONNECT SplitCLK_4_113_AND2T_18_n18(net143_c1,net143);
INTERCONNECT SplitCLK_4_113_OR2T_20_n20(net144_c1,net144);
INTERCONNECT SplitCLK_4_112_SplitCLK_6_108(net145_c1,net145);
INTERCONNECT SplitCLK_4_112_SplitCLK_4_111(net146_c1,net146);
INTERCONNECT SplitCLK_4_111_SplitCLK_4_109(net147_c1,net147);
INTERCONNECT SplitCLK_4_111_SplitCLK_4_110(net148_c1,net148);
INTERCONNECT SplitCLK_4_110_XOR2T_16_n16(net149_c1,net149);
INTERCONNECT SplitCLK_4_110_DFFT_69__FPB_n159(net150_c1,net150);
INTERCONNECT SplitCLK_4_109_AND2T_23_n23(net151_c1,net151);
INTERCONNECT SplitCLK_4_109_DFFT_70__FPB_n160(net152_c1,net152);
INTERCONNECT SplitCLK_6_108_SplitCLK_4_106(net153_c1,net153);
INTERCONNECT SplitCLK_6_108_SplitCLK_0_107(net154_c1,net154);
INTERCONNECT SplitCLK_0_107_XOR2T_21_n21(net155_c1,net155);
INTERCONNECT SplitCLK_0_107_DFFT_50__FPB_n140(net156_c1,net156);
INTERCONNECT SplitCLK_4_106_AND2T_24_n24(net157_c1,net157);
INTERCONNECT SplitCLK_4_106_OR2T_44_n44(net158_c1,net158);
INTERCONNECT SplitCLK_6_105_SplitCLK_4_98(net159_c1,net159);
INTERCONNECT SplitCLK_6_105_SplitCLK_2_104(net160_c1,net160);
INTERCONNECT SplitCLK_2_104_SplitCLK_2_101(net161_c1,net161);
INTERCONNECT SplitCLK_2_104_SplitCLK_4_103(net162_c1,net162);
INTERCONNECT SplitCLK_4_103_SplitCLK_2_123(net163_c1,net163);
INTERCONNECT SplitCLK_4_103_SplitCLK_4_102(net164_c1,net164);
INTERCONNECT SplitCLK_4_102_AND2T_25_n25(net165_c1,net165);
INTERCONNECT SplitCLK_4_102_OR2T_27_n27(net166_c1,net166);
INTERCONNECT SplitCLK_2_101_SplitCLK_4_99(net167_c1,net167);
INTERCONNECT SplitCLK_2_101_SplitCLK_4_100(net168_c1,net168);
INTERCONNECT SplitCLK_4_100_XOR2T_15_n15(net169_c1,net169);
INTERCONNECT SplitCLK_4_100_AND2T_19_n19(net170_c1,net170);
INTERCONNECT SplitCLK_4_99_AND2T_33_n33(net171_c1,net171);
INTERCONNECT SplitCLK_4_99_DFFT_58__FPB_n148(net172_c1,net172);
INTERCONNECT SplitCLK_4_98_SplitCLK_4_94(net173_c1,net173);
INTERCONNECT SplitCLK_4_98_SplitCLK_4_97(net174_c1,net174);
INTERCONNECT SplitCLK_4_97_SplitCLK_4_95(net175_c1,net175);
INTERCONNECT SplitCLK_4_97_SplitCLK_4_96(net176_c1,net176);
INTERCONNECT SplitCLK_4_96_AND2T_41_n41(net177_c1,net177);
INTERCONNECT SplitCLK_4_96_OR2T_35_n35(net178_c1,net178);
INTERCONNECT SplitCLK_4_95_DFFT_49__FPB_n139(net179_c1,net179);
INTERCONNECT SplitCLK_4_95_DFFT_59__FPB_n149(net180_c1,net180);
INTERCONNECT SplitCLK_4_94_SplitCLK_4_92(net181_c1,net181);
INTERCONNECT SplitCLK_4_94_SplitCLK_4_93(net182_c1,net182);
INTERCONNECT SplitCLK_4_93_AND2T_26_n26(net183_c1,net183);
INTERCONNECT SplitCLK_4_93_OR2T_43_n43(net184_c1,net184);
INTERCONNECT SplitCLK_4_92_XOR2T_17_n17(net185_c1,net185);
INTERCONNECT SplitCLK_4_92_DFFT_66__FPB_n156(net186_c1,net186);
INTERCONNECT SplitCLK_0_91_SplitCLK_2_76(net187_c1,net187);
INTERCONNECT SplitCLK_0_91_SplitCLK_4_90(net188_c1,net188);
INTERCONNECT SplitCLK_4_90_SplitCLK_0_83(net189_c1,net189);
INTERCONNECT SplitCLK_4_90_SplitCLK_4_89(net190_c1,net190);
INTERCONNECT SplitCLK_4_89_SplitCLK_6_86(net191_c1,net191);
INTERCONNECT SplitCLK_4_89_SplitCLK_4_88(net192_c1,net192);
INTERCONNECT SplitCLK_4_88_SplitCLK_2_121(net193_c1,net193);
INTERCONNECT SplitCLK_4_88_SplitCLK_4_87(net194_c1,net194);
INTERCONNECT SplitCLK_4_87_DFFT_74_sum1(net195_c1,net195);
INTERCONNECT SplitCLK_4_87_DFFT_71__FPB_n161(net196_c1,net196);
INTERCONNECT SplitCLK_6_86_SplitCLK_4_84(net197_c1,net197);
INTERCONNECT SplitCLK_6_86_SplitCLK_4_85(net198_c1,net198);
INTERCONNECT SplitCLK_4_85_AND2T_39_n39(net199_c1,net199);
INTERCONNECT SplitCLK_4_85_OR2T_45_cout(net200_c1,net200);
INTERCONNECT SplitCLK_4_84_DFFT_64__FPB_n154(net201_c1,net201);
INTERCONNECT SplitCLK_4_84_DFFT_68__FPB_n158(net202_c1,net202);
INTERCONNECT SplitCLK_0_83_SplitCLK_4_79(net203_c1,net203);
INTERCONNECT SplitCLK_0_83_SplitCLK_4_82(net204_c1,net204);
INTERCONNECT SplitCLK_4_82_SplitCLK_4_80(net205_c1,net205);
INTERCONNECT SplitCLK_4_82_SplitCLK_4_81(net206_c1,net206);
INTERCONNECT SplitCLK_4_81_AND2T_40_n40(net207_c1,net207);
INTERCONNECT SplitCLK_4_81_DFFT_73__FPB_n163(net208_c1,net208);
INTERCONNECT SplitCLK_4_80_OR2T_28_n28(net209_c1,net209);
INTERCONNECT SplitCLK_4_80_DFFT_75_sum2(net210_c1,net210);
INTERCONNECT SplitCLK_4_79_SplitCLK_4_77(net211_c1,net211);
INTERCONNECT SplitCLK_4_79_SplitCLK_4_78(net212_c1,net212);
INTERCONNECT SplitCLK_4_78_DFFT_55__FPB_n145(net213_c1,net213);
INTERCONNECT SplitCLK_4_78_DFFT_56__FPB_n146(net214_c1,net214);
INTERCONNECT SplitCLK_4_77_XOR2T_29_n29(net215_c1,net215);
INTERCONNECT SplitCLK_4_77_DFFT_65__FPB_n155(net216_c1,net216);
INTERCONNECT SplitCLK_2_76_SplitCLK_0_68(net217_c1,net217);
INTERCONNECT SplitCLK_2_76_SplitCLK_6_75(net218_c1,net218);
INTERCONNECT SplitCLK_6_75_SplitCLK_6_71(net219_c1,net219);
INTERCONNECT SplitCLK_6_75_SplitCLK_2_74(net220_c1,net220);
INTERCONNECT SplitCLK_2_74_SplitCLK_4_72(net221_c1,net221);
INTERCONNECT SplitCLK_2_74_SplitCLK_4_73(net222_c1,net222);
INTERCONNECT SplitCLK_4_73_AND2T_31_n31(net223_c1,net223);
INTERCONNECT SplitCLK_4_73_DFFT_67__FPB_n157(net224_c1,net224);
INTERCONNECT SplitCLK_4_72_AND2T_32_n32(net225_c1,net225);
INTERCONNECT SplitCLK_4_72_DFFT_57__FPB_n147(net226_c1,net226);
INTERCONNECT SplitCLK_6_71_SplitCLK_4_69(net227_c1,net227);
INTERCONNECT SplitCLK_6_71_SplitCLK_4_70(net228_c1,net228);
INTERCONNECT SplitCLK_4_70_XOR2T_22_n22(net229_c1,net229);
INTERCONNECT SplitCLK_4_70_AND2T_42_n42(net230_c1,net230);
INTERCONNECT SplitCLK_4_69_AND2T_34_n34(net231_c1,net231);
INTERCONNECT SplitCLK_4_69_AND2T_38_n38(net232_c1,net232);
INTERCONNECT SplitCLK_0_68_SplitCLK_6_64(net233_c1,net233);
INTERCONNECT SplitCLK_0_68_SplitCLK_4_67(net234_c1,net234);
INTERCONNECT SplitCLK_4_67_SplitCLK_4_65(net235_c1,net235);
INTERCONNECT SplitCLK_4_67_SplitCLK_4_66(net236_c1,net236);
INTERCONNECT SplitCLK_4_66_DFFT_61__FPB_n151(net237_c1,net237);
INTERCONNECT SplitCLK_4_66_DFFT_54__FPB_n144(net238_c1,net238);
INTERCONNECT SplitCLK_4_65_XOR2T_37_sum3(net239_c1,net239);
INTERCONNECT SplitCLK_4_65_OR2T_36_n36(net240_c1,net240);
INTERCONNECT SplitCLK_6_64_SplitCLK_4_62(net241_c1,net241);
INTERCONNECT SplitCLK_6_64_SplitCLK_4_63(net242_c1,net242);
INTERCONNECT SplitCLK_4_63_DFFT_60__FPB_n150(net243_c1,net243);
INTERCONNECT SplitCLK_4_63_DFFT_62__FPB_n152(net244_c1,net244);
INTERCONNECT SplitCLK_4_62_XOR2T_30_n30(net245_c1,net245);
INTERCONNECT SplitCLK_4_62_DFFT_63__FPB_n153(net246_c1,net246);
INTERCONNECT GCLK_Pad_SplitCLK_0_124(GCLK_Pad,net247);

endmodule
