`timescale 1ps / 1fs
module tb;
	reg GCLK_Pad;
	reg input1_Pad;
	reg input2_Pad;
	reg reset_Pad;
	wire state_obs0_Pad;
	wire state_obs1_Pad;
	wire output1_Pad;
	fsm1_route topLevel(.GCLK_Pad(GCLK_Pad), .input1_Pad(input1_Pad), .input2_Pad(input2_Pad), .reset_Pad(reset_Pad), .state_obs0_Pad(state_obs0_Pad), .state_obs1_Pad(state_obs1_Pad), .output1_Pad(output1_Pad));
	initial begin
		$dumpfile("fsm1_route.vcd");
		$dumpvars(0,tb);
		$sdf_annotate("fsm1_route_qVsim.sdf");
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#40;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd1;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd1;
		input2_Pad = 1'd1;
		reset_Pad = 1'd0;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd1;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd0;
		input2_Pad = 1'd1;
		reset_Pad = 1'd0;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd0;
		input2_Pad = 1'd1;
		reset_Pad = 1'd0;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd1;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd0;
		input2_Pad = 1'd1;
		reset_Pad = 1'd0;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd1;
		input2_Pad = 1'd1;
		reset_Pad = 1'd0;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd0;
		input2_Pad = 1'd1;
		reset_Pad = 1'd0;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd1;
		#2;
		input1_Pad = 1'd0;
		input2_Pad = 1'd0;
		reset_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#10 $finish;
	end
endmodule
