module fsm1_route(
input GCLK_Pad,
input input1_Pad,
input input2_Pad,
input reset_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output output1_Pad);

wire net0_c1;
wire state_obs0_Pad;
wire net1_c1;
wire state_obs1_Pad;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire reset_Pad;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire input1_Pad;
wire net137;
wire input2_Pad;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire output1_Pad;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire GCLK_Pad;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;

DFFT DFFT_99__FPB_n291(net287,net174,net181_c1);
SPLITT Split_162_state_obs0(net127,net204_c1,net0_c1);
XOR2T XOR2T_55_n70(net333,net38,net149,net29_c1);
SPLITT Split_157_output1(net133,net139_c1,net206_c1);
NOTT NOTT_8_n23(net349,net94,net4_c1);
NOTT NOTT_9_n24(net259,net101,net7_c1);
AND2T AND2T_10_n25(net361,net102,net178,net10_c1);
AND2T AND2T_20_n35(net399,net57,net162,net17_c1);
AND2T AND2T_21_n36(net317,net17,net13,net22_c1);
AND2T AND2T_30_n45(net403,net115,net72,net26_c1);
AND2T AND2T_22_n37(net222,net130,net173,net27_c1);
AND2T AND2T_15_n30(net331,net100,net121,net2_c1);
AND2T AND2T_23_n38(net303,net80,net177,net33_c1);
AND2T AND2T_16_n31(net363,net110,net113,net3_c1);
AND2T AND2T_40_n55(net251,net31,net71,net36_c1);
AND2T AND2T_32_n47(net429,net32,net169,net37_c1);
AND2T AND2T_24_n39(net357,net79,net183,net38_c1);
AND2T AND2T_17_n32(net239,net114,net14,net6_c1);
AND2T AND2T_41_n56(net313,net103,net194,net41_c1);
AND2T AND2T_26_n41(net221,net449,net161,net8_c1);
AND2T AND2T_50_n65(net220,net106,net105,net43_c1);
AND2T AND2T_35_n50(net277,net66,net45,net11_c1);
AND2T AND2T_43_n58(net219,net44,net200,net47_c1);
AND2T AND2T_36_n51(net278,net11,net42,net15_c1);
AND2T AND2T_29_n44(net237,net16,net187,net21_c1);
AND2T AND2T_53_n68(net415,net48,net156,net50_c1);
AND2T AND2T_46_n61(net293,net19,net150,net24_c1);
AND2T AND2T_38_n53(net383,net20,net201,net25_c1);
AND2T AND2T_54_n69(net411,net29,net159,net51_c1);
AND2T AND2T_56_n71(net417,net51,net151,net34_c1);
AND2T AND2T_48_n63(net439,net30,net152,net35_c1);
AND2T AND2T_57_n72(net245,net84,net153,net39_c1);
AND2T AND2T_49_n64(net425,net69,net88,net40_c1);
OR2T OR2T_11_n26(net233,net109,net158,net14_c1);
OR2T OR2T_12_n27(net371,net58,net160,net18_c1);
OR2T OR2T_31_n46(net218,net26,net89,net32_c1);
OR2T OR2T_25_n40(net249,net129,net191,net5_c1);
OR2T OR2T_33_n48(net271,net86,net176,net42_c1);
OR2T OR2T_42_n57(net319,net131,net199,net44_c1);
OR2T OR2T_34_n49(net275,net125,net182,net45_c1);
OR2T OR2T_27_n42(net265,net8,net27,net12_c1);
OR2T OR2T_19_n34(net358,net122,net99,net13_c1);
OR2T OR2T_51_n66(net404,net43,net63,net46_c1);
OR2T OR2T_28_n43(net260,net12,net165,net16_c1);
OR2T OR2T_52_n67(net437,net46,net154,net48_c1);
OR2T OR2T_44_n59(net294,net47,net41,net49_c1);
OR2T OR2T_45_n60(net288,net49,net202,net19_c1);
OR2T OR2T_37_n52(net426,net37,net186,net20_c1);
OR2T OR2T_47_n62(net416,net97,net124,net30_c1);
OR2T OR2T_39_n54(net246,net67,net181,net31_c1);
NOTT NOTT_13_n28(net325,net134,net23_c1);
NOTT NOTT_14_n29(net327,net136,net28_c1);
NOTT NOTT_18_n33(net217,net112,net9_c1);
DFFT DFFT_100__FPB_n292(net314,net132,net184_c1);
DFFT DFFT_101__FPB_n293(net332,net448,net188_c1);
DFFT DFFT_110__FPB_n302(net389,net146,net148_c1);
DFFT DFFT_102__FPB_n294(net326,net188,net194_c1);
DFFT DFFT_111__FPB_n303(net291,net148,net150_c1);
DFFT DFFT_103__FPB_n295(net405,net87,net195_c1);
DFFT DFFT_120__FPB_n312(net445,net78,net151_c1);
DFFT DFFT_112__FPB_n304(net216,net53,net152_c1);
DFFT DFFT_104__FPB_n296(net406,net195,net199_c1);
DFFT DFFT_121__FPB_n313(net215,net60,net153_c1);
DFFT DFFT_113__FPB_n305(net438,net40,net154_c1);
DFFT DFFT_105__FPB_n297(net320,net77,net200_c1);
DFFT DFFT_114__FPB_n306(net446,net123,net155_c1);
DFFT DFFT_106__FPB_n298(net214,net36,net202_c1);
DFFT DFFT_115__FPB_n307(net443,net155,net156_c1);
DFFT DFFT_107__FPB_n299(net384,net96,net203_c1);
DFFT DFFT_108__FPB_n300(net387,net203,net145_c1);
DFFT DFFT_116__FPB_n308(net440,net83,net157_c1);
DFFT DFFT_109__FPB_n301(net390,net145,net146_c1);
DFFT DFFT_117__FPB_n309(net418,net157,net159_c1);
DFFT DFFT_118__FPB_n310(net305,net135,net147_c1);
DFFT DFFT_119__FPB_n311(net328,net147,net149_c1);
DFFT DFFT_60__FBL_n252(net304,net24,net142_c1);
DFFT DFFT_61__FBL_n253(net400,net164,net143_c1);
DFFT DFFT_62__FBL_n254(net306,net172,net144_c1);
DFFT DFFT_70__FPB_n262(net334,net91,net162_c1);
DFFT DFFT_71__FPB_n263(net351,net111,net163_c1);
DFFT DFFT_63__FPB_n255(net213,net50,net164_c1);
DFFT DFFT_80__FPB_n272(net345,net95,net166_c1);
DFFT DFFT_72__FPB_n264(net352,net163,net167_c1);
DFFT DFFT_64__FPB_n256(net412,net34,net168_c1);
DFFT DFFT_81__FPB_n273(net212,net166,net171_c1);
DFFT DFFT_73__FPB_n265(net372,net167,net173_c1);
DFFT DFFT_65__FPB_n257(net299,net168,net172_c1);
DFFT DFFT_58__FBL_n250(net238,net21,net140_c1);
DFFT DFFT_90__FPB_n282(net252,net170,net176_c1);
DFFT DFFT_82__FPB_n274(net263,net171,net175_c1);
DFFT DFFT_74__FPB_n266(net300,net93,net177_c1);
DFFT DFFT_66__FPB_n258(net362,net70,net178_c1);
DFFT DFFT_59__FBL_n251(net318,net25,net141_c1);
SPLITT Split_122_n314(net137,net54_c1,net98_c1);
SPLITT Split_130_n322(net7,net56_c1,net99_c1);
SPLITT Split_123_n315(net98,net59_c1,net101_c1);
SPLITT Split_131_n323(net56,net58_c1,net102_c1);
SPLITT Split_124_n316(net54,net60_c1,net104_c1);
SPLITT Split_132_n324(net10,net61_c1,net105_c1);
SPLITT Split_140_n332(net2,net62_c1,net106_c1);
SPLITT Split_125_n317(net138,net65_c1,net108_c1);
SPLITT Split_133_n325(net61,net67_c1,net109_c1);
SPLITT Split_141_n333(net62,net66_c1,net110_c1);
SPLITT Split_126_n318(net65,net70_c1,net112_c1);
SPLITT Split_134_n326(net18,net72_c1,net113_c1);
SPLITT Split_142_n334(net3,net71_c1,net114_c1);
SPLITT Split_150_n342(net107,net69_c1,net115_c1);
SPLITT Split_127_n319(net4,net75_c1,net117_c1);
SPLITT Split_135_n327(net23,net74_c1,net118_c1);
SPLITT Split_143_n335(net9,net73_c1,net119_c1);
SPLITT Split_151_n343(net64,net77_c1,net120_c1);
SPLITT Split_128_n320(net117,net52_c1,net95_c1);
SPLITT Split_136_n328(net118,net80_c1,net121_c1);
SPLITT Split_144_n336(net119,net79_c1,net122_c1);
SPLITT Split_152_n344(net35,net78_c1,net123_c1);
SPLITT Split_129_n321(net75,net53_c1,net96_c1);
SPLITT Split_137_n329(net74,net83_c1,net124_c1);
SPLITT Split_145_n337(net73,net84_c1,net125_c1);
SPLITT Split_153_n345(net39,net82_c1,net126_c1);
SPLITT Split_161_n353(net142,net81_c1,net127_c1);
SPLITT Split_138_n330(net28,net55_c1,net97_c1);
SPLITT Split_146_n338(net22,net85_c1,net128_c1);
SPLITT Split_154_n346(net126,net86_c1,net129_c1);
SPLITT Split_139_n331(net55,net57_c1,net100_c1);
SPLITT Split_147_n339(net128,net89_c1,net130_c1);
SPLITT Split_155_n347(net82,net88_c1,net131_c1);
SPLITT Split_163_n355(net81,net87_c1,net132_c1);
SPLITT Split_148_n340(net85,net63_c1,net103_c1);
SPLITT Split_156_n348(net140,net90_c1,net133_c1);
SPLITT Split_164_n356(net143,net91_c1,net134_c1);
SPLITT Split_149_n341(net33,net64_c1,net107_c1);
SPLITT Split_165_n357(net144,net92_c1,net135_c1);
SPLITT Split_158_n350(net90,net68_c1,net111_c1);
SPLITT Split_166_n358(net92,net93_c1,net136_c1);
SPLITT Split_159_n351(net141,net76_c1,net116_c1);
DFFT DFFT_91__FPB_n283(net250,net104,net182_c1);
DFFT DFFT_83__FPB_n275(net264,net175,net179_c1);
DFFT DFFT_75__FPB_n267(net276,net59,net183_c1);
DFFT DFFT_67__FPB_n259(net211,net139,net180_c1);
DFFT DFFT_68__FPB_n260(net234,net180,net158_c1);
DFFT DFFT_92__FPB_n284(net364,net15,net186_c1);
DFFT DFFT_84__FPB_n276(net210,net179,net187_c1);
DFFT DFFT_76__FPB_n268(net266,net68,net185_c1);
DFFT DFFT_69__FPB_n261(net377,net108,net160_c1);
DFFT DFFT_93__FPB_n285(net350,net52,net189_c1);
DFFT DFFT_85__FPB_n277(net444,net205,net190_c1);
DFFT DFFT_77__FPB_n269(net346,net185,net191_c1);
DFFT DFFT_78__FPB_n270(net272,net120,net161_c1);
DFFT DFFT_94__FPB_n286(net375,net189,net192_c1);
DFFT DFFT_86__FPB_n278(net431,net190,net193_c1);
DFFT DFFT_79__FPB_n271(net240,net6,net165_c1);
DFFT DFFT_95__FPB_n287(net378,net192,net196_c1);
DFFT DFFT_87__FPB_n279(net432,net193,net197_c1);
DFFT DFFT_88__FPB_n280(net430,net197,net169_c1);
DFFT DFFT_96__FPB_n288(net376,net196,net198_c1);
DFFT DFFT_89__FPB_n281(net292,net116,net170_c1);
DFFT DFFT_97__FPB_n289(net388,net198,net201_c1);
SPLITT Split_160_state_obs1(net76,net205_c1,net1_c1);
DFFT DFFT_98__FPB_n290(net209,net204,net174_c1);
SPLITT SplitCLK_4_115(net441,net445_c1,net446_c1);
SPLITT SplitCLK_4_116(net442,net443_c1,net444_c1);
SPLITT SplitCLK_4_117(net433,net441_c1,net442_c1);
SPLITT SplitCLK_4_118(net435,net439_c1,net440_c1);
SPLITT SplitCLK_4_119(net436,net437_c1,net438_c1);
SPLITT SplitCLK_2_120(net434,net436_c1,net435_c1);
SPLITT SplitCLK_6_121(net419,net433_c1,net434_c1);
SPLITT SplitCLK_0_122(net427,net431_c1,net432_c1);
SPLITT SplitCLK_4_123(net428,net429_c1,net430_c1);
SPLITT SplitCLK_0_124(net421,net427_c1,net428_c1);
SPLITT SplitCLK_4_125(net424,net425_c1,net426_c1);
SPLITT SplitCLK_6_126(net422,net424_c1,net423_c1);
SPLITT SplitCLK_4_127(net420,net422_c1,net421_c1);
SPLITT SplitCLK_0_128(net391,net419_c1,net420_c1);
SPLITT SplitCLK_0_129(net413,net417_c1,net418_c1);
SPLITT SplitCLK_4_130(net414,net415_c1,net416_c1);
SPLITT SplitCLK_0_131(net407,net413_c1,net414_c1);
SPLITT SplitCLK_4_132(net410,net412_c1,net411_c1);
SPLITT SplitCLK_2_133(net408,net409_c1,net410_c1);
SPLITT SplitCLK_6_134(net393,net407_c1,net408_c1);
SPLITT SplitCLK_4_135(net401,net406_c1,net405_c1);
SPLITT SplitCLK_4_136(net402,net403_c1,net404_c1);
SPLITT SplitCLK_0_137(net395,net401_c1,net402_c1);
SPLITT SplitCLK_4_138(net398,net400_c1,net399_c1);
SPLITT SplitCLK_2_139(net396,net397_c1,net398_c1);
SPLITT SplitCLK_6_140(net394,net395_c1,net396_c1);
SPLITT SplitCLK_6_141(net392,net393_c1,net394_c1);
SPLITT SplitCLK_6_142(net335,net391_c1,net392_c1);
SPLITT SplitCLK_4_143(net385,net389_c1,net390_c1);
SPLITT SplitCLK_4_144(net386,net388_c1,net387_c1);
SPLITT SplitCLK_6_145(net379,net385_c1,net386_c1);
SPLITT SplitCLK_4_146(net382,net383_c1,net384_c1);
SPLITT SplitCLK_2_147(net380,net381_c1,net382_c1);
SPLITT SplitCLK_4_148(net365,net380_c1,net379_c1);
SPLITT SplitCLK_4_149(net373,net377_c1,net378_c1);
SPLITT SplitCLK_4_150(net374,net375_c1,net376_c1);
SPLITT SplitCLK_4_151(net367,net374_c1,net373_c1);
SPLITT SplitCLK_4_152(net370,net371_c1,net372_c1);
SPLITT SplitCLK_2_153(net368,net369_c1,net370_c1);
SPLITT SplitCLK_4_154(net366,net368_c1,net367_c1);
SPLITT SplitCLK_0_155(net337,net365_c1,net366_c1);
SPLITT SplitCLK_0_156(net359,net363_c1,net364_c1);
SPLITT SplitCLK_4_157(net360,net362_c1,net361_c1);
SPLITT SplitCLK_0_158(net353,net359_c1,net360_c1);
SPLITT SplitCLK_4_159(net356,net357_c1,net358_c1);
SPLITT SplitCLK_6_160(net354,net356_c1,net355_c1);
SPLITT SplitCLK_6_161(net339,net353_c1,net354_c1);
SPLITT SplitCLK_0_162(net347,net351_c1,net352_c1);
SPLITT SplitCLK_4_163(net348,net350_c1,net349_c1);
SPLITT SplitCLK_0_164(net341,net347_c1,net348_c1);
SPLITT SplitCLK_4_165(net344,net345_c1,net346_c1);
SPLITT SplitCLK_6_166(net342,net344_c1,net343_c1);
SPLITT SplitCLK_4_167(net340,net342_c1,net341_c1);
SPLITT SplitCLK_4_168(net338,net340_c1,net339_c1);
SPLITT SplitCLK_4_169(net336,net338_c1,net337_c1);
SPLITT SplitCLK_0_170(net207,net335_c1,net336_c1);
SPLITT SplitCLK_4_171(net329,net334_c1,net333_c1);
SPLITT SplitCLK_4_172(net330,net332_c1,net331_c1);
SPLITT SplitCLK_4_173(net321,net329_c1,net330_c1);
SPLITT SplitCLK_0_174(net323,net327_c1,net328_c1);
SPLITT SplitCLK_4_175(net324,net325_c1,net326_c1);
SPLITT SplitCLK_6_176(net322,net324_c1,net323_c1);
SPLITT SplitCLK_6_177(net307,net321_c1,net322_c1);
SPLITT SplitCLK_4_178(net315,net319_c1,net320_c1);
SPLITT SplitCLK_4_179(net316,net318_c1,net317_c1);
SPLITT SplitCLK_0_180(net309,net315_c1,net316_c1);
SPLITT SplitCLK_4_181(net312,net314_c1,net313_c1);
SPLITT SplitCLK_2_182(net310,net311_c1,net312_c1);
SPLITT SplitCLK_4_183(net308,net310_c1,net309_c1);
SPLITT SplitCLK_0_184(net279,net307_c1,net308_c1);
SPLITT SplitCLK_0_185(net301,net305_c1,net306_c1);
SPLITT SplitCLK_4_186(net302,net303_c1,net304_c1);
SPLITT SplitCLK_4_187(net295,net302_c1,net301_c1);
SPLITT SplitCLK_4_188(net298,net299_c1,net300_c1);
SPLITT SplitCLK_2_189(net296,net297_c1,net298_c1);
SPLITT SplitCLK_6_190(net281,net295_c1,net296_c1);
SPLITT SplitCLK_0_191(net289,net293_c1,net294_c1);
SPLITT SplitCLK_4_192(net290,net291_c1,net292_c1);
SPLITT SplitCLK_0_193(net283,net289_c1,net290_c1);
SPLITT SplitCLK_4_194(net286,net287_c1,net288_c1);
SPLITT SplitCLK_2_195(net284,net285_c1,net286_c1);
SPLITT SplitCLK_4_196(net282,net284_c1,net283_c1);
SPLITT SplitCLK_2_197(net280,net282_c1,net281_c1);
SPLITT SplitCLK_6_198(net223,net279_c1,net280_c1);
SPLITT SplitCLK_4_199(net273,net278_c1,net277_c1);
SPLITT SplitCLK_4_200(net274,net276_c1,net275_c1);
SPLITT SplitCLK_0_201(net267,net273_c1,net274_c1);
SPLITT SplitCLK_4_202(net270,net271_c1,net272_c1);
SPLITT SplitCLK_2_203(net268,net269_c1,net270_c1);
SPLITT SplitCLK_2_204(net253,net267_c1,net268_c1);
SPLITT SplitCLK_4_205(net261,net265_c1,net266_c1);
SPLITT SplitCLK_4_206(net262,net264_c1,net263_c1);
SPLITT SplitCLK_0_207(net255,net261_c1,net262_c1);
SPLITT SplitCLK_4_208(net258,net259_c1,net260_c1);
SPLITT SplitCLK_2_209(net256,net257_c1,net258_c1);
SPLITT SplitCLK_4_210(net254,net256_c1,net255_c1);
SPLITT SplitCLK_0_211(net225,net253_c1,net254_c1);
SPLITT SplitCLK_0_212(net247,net251_c1,net252_c1);
SPLITT SplitCLK_4_213(net248,net250_c1,net249_c1);
SPLITT SplitCLK_0_214(net241,net247_c1,net248_c1);
SPLITT SplitCLK_4_215(net244,net246_c1,net245_c1);
SPLITT SplitCLK_2_216(net242,net243_c1,net244_c1);
SPLITT SplitCLK_6_217(net227,net241_c1,net242_c1);
SPLITT SplitCLK_4_218(net235,net239_c1,net240_c1);
SPLITT SplitCLK_4_219(net236,net238_c1,net237_c1);
SPLITT SplitCLK_4_220(net229,net235_c1,net236_c1);
SPLITT SplitCLK_4_221(net232,net234_c1,net233_c1);
SPLITT SplitCLK_2_222(net230,net231_c1,net232_c1);
SPLITT SplitCLK_4_223(net228,net230_c1,net229_c1);
SPLITT SplitCLK_2_224(net226,net228_c1,net227_c1);
SPLITT SplitCLK_4_225(net224,net226_c1,net225_c1);
SPLITT SplitCLK_2_226(net208,net224_c1,net223_c1);
wire dummy0;
SPLITT SplitCLK_2_227(net369,net222_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_4_228(net269,net221_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_4_229(net397,net220_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_230(net311,net219_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_231(net423,net218_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_4_232(net355,net217_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_2_233(net381,net216_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_4_234(net243,net215_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_2_235(net285,net214_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_4_236(net409,net213_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_2_237(net343,net212_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_4_238(net231,net211_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_4_239(net257,net210_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_4_240(net297,net209_c1,dummy13);
SPLITT SplitCLK_0_241(net447,net207_c1,net208_c1);
wire dummy14;
SPLITT Split_HOLD_294(net184,dummy14,net448_c1);
wire dummy15;
SPLITT Split_HOLD_295(net5,dummy15,net449_c1);
INTERCONNECT Split_162_state_obs0_state_obs0_Pad(net0_c1,state_obs0_Pad);
INTERCONNECT Split_160_state_obs1_state_obs1_Pad(net1_c1,state_obs1_Pad);
INTERCONNECT AND2T_15_n30_Split_140_n332(net2_c1,net2);
INTERCONNECT AND2T_16_n31_Split_142_n334(net3_c1,net3);
INTERCONNECT NOTT_8_n23_Split_127_n319(net4_c1,net4);
INTERCONNECT OR2T_25_n40_Split_HOLD_295(net5_c1,net5);
INTERCONNECT AND2T_17_n32_DFFT_79__FPB_n271(net6_c1,net6);
INTERCONNECT NOTT_9_n24_Split_130_n322(net7_c1,net7);
INTERCONNECT AND2T_26_n41_OR2T_27_n42(net8_c1,net8);
INTERCONNECT NOTT_18_n33_Split_143_n335(net9_c1,net9);
INTERCONNECT AND2T_10_n25_Split_132_n324(net10_c1,net10);
INTERCONNECT AND2T_35_n50_AND2T_36_n51(net11_c1,net11);
INTERCONNECT OR2T_27_n42_OR2T_28_n43(net12_c1,net12);
INTERCONNECT OR2T_19_n34_AND2T_21_n36(net13_c1,net13);
INTERCONNECT OR2T_11_n26_AND2T_17_n32(net14_c1,net14);
INTERCONNECT AND2T_36_n51_DFFT_92__FPB_n284(net15_c1,net15);
INTERCONNECT OR2T_28_n43_AND2T_29_n44(net16_c1,net16);
INTERCONNECT AND2T_20_n35_AND2T_21_n36(net17_c1,net17);
INTERCONNECT OR2T_12_n27_Split_134_n326(net18_c1,net18);
INTERCONNECT OR2T_45_n60_AND2T_46_n61(net19_c1,net19);
INTERCONNECT OR2T_37_n52_AND2T_38_n53(net20_c1,net20);
INTERCONNECT AND2T_29_n44_DFFT_58__FBL_n250(net21_c1,net21);
INTERCONNECT AND2T_21_n36_Split_146_n338(net22_c1,net22);
INTERCONNECT NOTT_13_n28_Split_135_n327(net23_c1,net23);
INTERCONNECT AND2T_46_n61_DFFT_60__FBL_n252(net24_c1,net24);
INTERCONNECT AND2T_38_n53_DFFT_59__FBL_n251(net25_c1,net25);
INTERCONNECT AND2T_30_n45_OR2T_31_n46(net26_c1,net26);
INTERCONNECT AND2T_22_n37_OR2T_27_n42(net27_c1,net27);
INTERCONNECT NOTT_14_n29_Split_138_n330(net28_c1,net28);
INTERCONNECT XOR2T_55_n70_AND2T_54_n69(net29_c1,net29);
INTERCONNECT OR2T_47_n62_AND2T_48_n63(net30_c1,net30);
INTERCONNECT OR2T_39_n54_AND2T_40_n55(net31_c1,net31);
INTERCONNECT OR2T_31_n46_AND2T_32_n47(net32_c1,net32);
INTERCONNECT AND2T_23_n38_Split_149_n341(net33_c1,net33);
INTERCONNECT AND2T_56_n71_DFFT_64__FPB_n256(net34_c1,net34);
INTERCONNECT AND2T_48_n63_Split_152_n344(net35_c1,net35);
INTERCONNECT AND2T_40_n55_DFFT_106__FPB_n298(net36_c1,net36);
INTERCONNECT AND2T_32_n47_OR2T_37_n52(net37_c1,net37);
INTERCONNECT AND2T_24_n39_XOR2T_55_n70(net38_c1,net38);
INTERCONNECT AND2T_57_n72_Split_153_n345(net39_c1,net39);
INTERCONNECT AND2T_49_n64_DFFT_113__FPB_n305(net40_c1,net40);
INTERCONNECT AND2T_41_n56_OR2T_44_n59(net41_c1,net41);
INTERCONNECT OR2T_33_n48_AND2T_36_n51(net42_c1,net42);
INTERCONNECT AND2T_50_n65_OR2T_51_n66(net43_c1,net43);
INTERCONNECT OR2T_42_n57_AND2T_43_n58(net44_c1,net44);
INTERCONNECT OR2T_34_n49_AND2T_35_n50(net45_c1,net45);
INTERCONNECT OR2T_51_n66_OR2T_52_n67(net46_c1,net46);
INTERCONNECT AND2T_43_n58_OR2T_44_n59(net47_c1,net47);
INTERCONNECT OR2T_52_n67_AND2T_53_n68(net48_c1,net48);
INTERCONNECT OR2T_44_n59_OR2T_45_n60(net49_c1,net49);
INTERCONNECT AND2T_53_n68_DFFT_63__FPB_n255(net50_c1,net50);
INTERCONNECT AND2T_54_n69_AND2T_56_n71(net51_c1,net51);
INTERCONNECT Split_128_n320_DFFT_93__FPB_n285(net52_c1,net52);
INTERCONNECT Split_129_n321_DFFT_112__FPB_n304(net53_c1,net53);
INTERCONNECT Split_122_n314_Split_124_n316(net54_c1,net54);
INTERCONNECT Split_138_n330_Split_139_n331(net55_c1,net55);
INTERCONNECT Split_130_n322_Split_131_n323(net56_c1,net56);
INTERCONNECT Split_139_n331_AND2T_20_n35(net57_c1,net57);
INTERCONNECT Split_131_n323_OR2T_12_n27(net58_c1,net58);
INTERCONNECT Split_123_n315_DFFT_75__FPB_n267(net59_c1,net59);
INTERCONNECT Split_124_n316_DFFT_121__FPB_n313(net60_c1,net60);
INTERCONNECT Split_132_n324_Split_133_n325(net61_c1,net61);
INTERCONNECT Split_140_n332_Split_141_n333(net62_c1,net62);
INTERCONNECT Split_148_n340_OR2T_51_n66(net63_c1,net63);
INTERCONNECT Split_149_n341_Split_151_n343(net64_c1,net64);
INTERCONNECT Split_125_n317_Split_126_n318(net65_c1,net65);
INTERCONNECT Split_141_n333_AND2T_35_n50(net66_c1,net66);
INTERCONNECT Split_133_n325_OR2T_39_n54(net67_c1,net67);
INTERCONNECT Split_158_n350_DFFT_76__FPB_n268(net68_c1,net68);
INTERCONNECT Split_150_n342_AND2T_49_n64(net69_c1,net69);
INTERCONNECT Split_126_n318_DFFT_66__FPB_n258(net70_c1,net70);
INTERCONNECT Split_142_n334_AND2T_40_n55(net71_c1,net71);
INTERCONNECT Split_134_n326_AND2T_30_n45(net72_c1,net72);
INTERCONNECT Split_143_n335_Split_145_n337(net73_c1,net73);
INTERCONNECT Split_135_n327_Split_137_n329(net74_c1,net74);
INTERCONNECT Split_127_n319_Split_129_n321(net75_c1,net75);
INTERCONNECT Split_159_n351_Split_160_state_obs1(net76_c1,net76);
INTERCONNECT Split_151_n343_DFFT_105__FPB_n297(net77_c1,net77);
INTERCONNECT Split_152_n344_DFFT_120__FPB_n312(net78_c1,net78);
INTERCONNECT Split_144_n336_AND2T_24_n39(net79_c1,net79);
INTERCONNECT Split_136_n328_AND2T_23_n38(net80_c1,net80);
INTERCONNECT Split_161_n353_Split_163_n355(net81_c1,net81);
INTERCONNECT Split_153_n345_Split_155_n347(net82_c1,net82);
INTERCONNECT Split_137_n329_DFFT_116__FPB_n308(net83_c1,net83);
INTERCONNECT Split_145_n337_AND2T_57_n72(net84_c1,net84);
INTERCONNECT Split_146_n338_Split_148_n340(net85_c1,net85);
INTERCONNECT Split_154_n346_OR2T_33_n48(net86_c1,net86);
INTERCONNECT Split_163_n355_DFFT_103__FPB_n295(net87_c1,net87);
INTERCONNECT Split_155_n347_AND2T_49_n64(net88_c1,net88);
INTERCONNECT Split_147_n339_OR2T_31_n46(net89_c1,net89);
INTERCONNECT Split_156_n348_Split_158_n350(net90_c1,net90);
INTERCONNECT Split_164_n356_DFFT_70__FPB_n262(net91_c1,net91);
INTERCONNECT Split_165_n357_Split_166_n358(net92_c1,net92);
INTERCONNECT Split_166_n358_DFFT_74__FPB_n266(net93_c1,net93);
INTERCONNECT reset_Pad_NOTT_8_n23(reset_Pad,net94);
INTERCONNECT Split_128_n320_DFFT_80__FPB_n272(net95_c1,net95);
INTERCONNECT Split_129_n321_DFFT_107__FPB_n299(net96_c1,net96);
INTERCONNECT Split_138_n330_OR2T_47_n62(net97_c1,net97);
INTERCONNECT Split_122_n314_Split_123_n315(net98_c1,net98);
INTERCONNECT Split_130_n322_OR2T_19_n34(net99_c1,net99);
INTERCONNECT Split_139_n331_AND2T_15_n30(net100_c1,net100);
INTERCONNECT Split_123_n315_NOTT_9_n24(net101_c1,net101);
INTERCONNECT Split_131_n323_AND2T_10_n25(net102_c1,net102);
INTERCONNECT Split_148_n340_AND2T_41_n56(net103_c1,net103);
INTERCONNECT Split_124_n316_DFFT_91__FPB_n283(net104_c1,net104);
INTERCONNECT Split_132_n324_AND2T_50_n65(net105_c1,net105);
INTERCONNECT Split_140_n332_AND2T_50_n65(net106_c1,net106);
INTERCONNECT Split_149_n341_Split_150_n342(net107_c1,net107);
INTERCONNECT Split_125_n317_DFFT_69__FPB_n261(net108_c1,net108);
INTERCONNECT Split_133_n325_OR2T_11_n26(net109_c1,net109);
INTERCONNECT Split_141_n333_AND2T_16_n31(net110_c1,net110);
INTERCONNECT Split_158_n350_DFFT_71__FPB_n263(net111_c1,net111);
INTERCONNECT Split_126_n318_NOTT_18_n33(net112_c1,net112);
INTERCONNECT Split_134_n326_AND2T_16_n31(net113_c1,net113);
INTERCONNECT Split_142_n334_AND2T_17_n32(net114_c1,net114);
INTERCONNECT Split_150_n342_AND2T_30_n45(net115_c1,net115);
INTERCONNECT Split_159_n351_DFFT_89__FPB_n281(net116_c1,net116);
INTERCONNECT Split_127_n319_Split_128_n320(net117_c1,net117);
INTERCONNECT Split_135_n327_Split_136_n328(net118_c1,net118);
INTERCONNECT Split_143_n335_Split_144_n336(net119_c1,net119);
INTERCONNECT Split_151_n343_DFFT_78__FPB_n270(net120_c1,net120);
INTERCONNECT Split_136_n328_AND2T_15_n30(net121_c1,net121);
INTERCONNECT Split_144_n336_OR2T_19_n34(net122_c1,net122);
INTERCONNECT Split_152_n344_DFFT_114__FPB_n306(net123_c1,net123);
INTERCONNECT Split_137_n329_OR2T_47_n62(net124_c1,net124);
INTERCONNECT Split_145_n337_OR2T_34_n49(net125_c1,net125);
INTERCONNECT Split_153_n345_Split_154_n346(net126_c1,net126);
INTERCONNECT Split_161_n353_Split_162_state_obs0(net127_c1,net127);
INTERCONNECT Split_146_n338_Split_147_n339(net128_c1,net128);
INTERCONNECT Split_154_n346_OR2T_25_n40(net129_c1,net129);
INTERCONNECT Split_147_n339_AND2T_22_n37(net130_c1,net130);
INTERCONNECT Split_155_n347_OR2T_42_n57(net131_c1,net131);
INTERCONNECT Split_163_n355_DFFT_100__FPB_n292(net132_c1,net132);
INTERCONNECT Split_156_n348_Split_157_output1(net133_c1,net133);
INTERCONNECT Split_164_n356_NOTT_13_n28(net134_c1,net134);
INTERCONNECT Split_165_n357_DFFT_118__FPB_n310(net135_c1,net135);
INTERCONNECT Split_166_n358_NOTT_14_n29(net136_c1,net136);
INTERCONNECT input1_Pad_Split_122_n314(input1_Pad,net137);
INTERCONNECT input2_Pad_Split_125_n317(input2_Pad,net138);
INTERCONNECT Split_157_output1_DFFT_67__FPB_n259(net139_c1,net139);
INTERCONNECT DFFT_58__FBL_n250_Split_156_n348(net140_c1,net140);
INTERCONNECT DFFT_59__FBL_n251_Split_159_n351(net141_c1,net141);
INTERCONNECT DFFT_60__FBL_n252_Split_161_n353(net142_c1,net142);
INTERCONNECT DFFT_61__FBL_n253_Split_164_n356(net143_c1,net143);
INTERCONNECT DFFT_62__FBL_n254_Split_165_n357(net144_c1,net144);
INTERCONNECT DFFT_108__FPB_n300_DFFT_109__FPB_n301(net145_c1,net145);
INTERCONNECT DFFT_109__FPB_n301_DFFT_110__FPB_n302(net146_c1,net146);
INTERCONNECT DFFT_118__FPB_n310_DFFT_119__FPB_n311(net147_c1,net147);
INTERCONNECT DFFT_110__FPB_n302_DFFT_111__FPB_n303(net148_c1,net148);
INTERCONNECT DFFT_119__FPB_n311_XOR2T_55_n70(net149_c1,net149);
INTERCONNECT DFFT_111__FPB_n303_AND2T_46_n61(net150_c1,net150);
INTERCONNECT DFFT_120__FPB_n312_AND2T_56_n71(net151_c1,net151);
INTERCONNECT DFFT_112__FPB_n304_AND2T_48_n63(net152_c1,net152);
INTERCONNECT DFFT_121__FPB_n313_AND2T_57_n72(net153_c1,net153);
INTERCONNECT DFFT_113__FPB_n305_OR2T_52_n67(net154_c1,net154);
INTERCONNECT DFFT_114__FPB_n306_DFFT_115__FPB_n307(net155_c1,net155);
INTERCONNECT DFFT_115__FPB_n307_AND2T_53_n68(net156_c1,net156);
INTERCONNECT DFFT_116__FPB_n308_DFFT_117__FPB_n309(net157_c1,net157);
INTERCONNECT DFFT_68__FPB_n260_OR2T_11_n26(net158_c1,net158);
INTERCONNECT DFFT_117__FPB_n309_AND2T_54_n69(net159_c1,net159);
INTERCONNECT DFFT_69__FPB_n261_OR2T_12_n27(net160_c1,net160);
INTERCONNECT DFFT_78__FPB_n270_AND2T_26_n41(net161_c1,net161);
INTERCONNECT DFFT_70__FPB_n262_AND2T_20_n35(net162_c1,net162);
INTERCONNECT DFFT_71__FPB_n263_DFFT_72__FPB_n264(net163_c1,net163);
INTERCONNECT DFFT_63__FPB_n255_DFFT_61__FBL_n253(net164_c1,net164);
INTERCONNECT DFFT_79__FPB_n271_OR2T_28_n43(net165_c1,net165);
INTERCONNECT DFFT_80__FPB_n272_DFFT_81__FPB_n273(net166_c1,net166);
INTERCONNECT DFFT_72__FPB_n264_DFFT_73__FPB_n265(net167_c1,net167);
INTERCONNECT DFFT_64__FPB_n256_DFFT_65__FPB_n257(net168_c1,net168);
INTERCONNECT DFFT_88__FPB_n280_AND2T_32_n47(net169_c1,net169);
INTERCONNECT DFFT_89__FPB_n281_DFFT_90__FPB_n282(net170_c1,net170);
INTERCONNECT DFFT_81__FPB_n273_DFFT_82__FPB_n274(net171_c1,net171);
INTERCONNECT DFFT_65__FPB_n257_DFFT_62__FBL_n254(net172_c1,net172);
INTERCONNECT DFFT_73__FPB_n265_AND2T_22_n37(net173_c1,net173);
INTERCONNECT DFFT_98__FPB_n290_DFFT_99__FPB_n291(net174_c1,net174);
INTERCONNECT DFFT_82__FPB_n274_DFFT_83__FPB_n275(net175_c1,net175);
INTERCONNECT DFFT_90__FPB_n282_OR2T_33_n48(net176_c1,net176);
INTERCONNECT DFFT_74__FPB_n266_AND2T_23_n38(net177_c1,net177);
INTERCONNECT DFFT_66__FPB_n258_AND2T_10_n25(net178_c1,net178);
INTERCONNECT DFFT_83__FPB_n275_DFFT_84__FPB_n276(net179_c1,net179);
INTERCONNECT DFFT_67__FPB_n259_DFFT_68__FPB_n260(net180_c1,net180);
INTERCONNECT DFFT_99__FPB_n291_OR2T_39_n54(net181_c1,net181);
INTERCONNECT DFFT_91__FPB_n283_OR2T_34_n49(net182_c1,net182);
INTERCONNECT DFFT_75__FPB_n267_AND2T_24_n39(net183_c1,net183);
INTERCONNECT DFFT_100__FPB_n292_Split_HOLD_294(net184_c1,net184);
INTERCONNECT DFFT_76__FPB_n268_DFFT_77__FPB_n269(net185_c1,net185);
INTERCONNECT DFFT_92__FPB_n284_OR2T_37_n52(net186_c1,net186);
INTERCONNECT DFFT_84__FPB_n276_AND2T_29_n44(net187_c1,net187);
INTERCONNECT DFFT_101__FPB_n293_DFFT_102__FPB_n294(net188_c1,net188);
INTERCONNECT DFFT_93__FPB_n285_DFFT_94__FPB_n286(net189_c1,net189);
INTERCONNECT DFFT_85__FPB_n277_DFFT_86__FPB_n278(net190_c1,net190);
INTERCONNECT DFFT_77__FPB_n269_OR2T_25_n40(net191_c1,net191);
INTERCONNECT DFFT_94__FPB_n286_DFFT_95__FPB_n287(net192_c1,net192);
INTERCONNECT DFFT_86__FPB_n278_DFFT_87__FPB_n279(net193_c1,net193);
INTERCONNECT DFFT_102__FPB_n294_AND2T_41_n56(net194_c1,net194);
INTERCONNECT DFFT_103__FPB_n295_DFFT_104__FPB_n296(net195_c1,net195);
INTERCONNECT DFFT_95__FPB_n287_DFFT_96__FPB_n288(net196_c1,net196);
INTERCONNECT DFFT_87__FPB_n279_DFFT_88__FPB_n280(net197_c1,net197);
INTERCONNECT DFFT_96__FPB_n288_DFFT_97__FPB_n289(net198_c1,net198);
INTERCONNECT DFFT_104__FPB_n296_OR2T_42_n57(net199_c1,net199);
INTERCONNECT DFFT_105__FPB_n297_AND2T_43_n58(net200_c1,net200);
INTERCONNECT DFFT_97__FPB_n289_AND2T_38_n53(net201_c1,net201);
INTERCONNECT DFFT_106__FPB_n298_OR2T_45_n60(net202_c1,net202);
INTERCONNECT DFFT_107__FPB_n299_DFFT_108__FPB_n300(net203_c1,net203);
INTERCONNECT Split_162_state_obs0_DFFT_98__FPB_n290(net204_c1,net204);
INTERCONNECT Split_160_state_obs1_DFFT_85__FPB_n277(net205_c1,net205);
INTERCONNECT Split_157_output1_output1_Pad(net206_c1,output1_Pad);
INTERCONNECT SplitCLK_0_241_SplitCLK_0_170(net207_c1,net207);
INTERCONNECT SplitCLK_0_241_SplitCLK_2_226(net208_c1,net208);
INTERCONNECT SplitCLK_4_240_DFFT_98__FPB_n290(net209_c1,net209);
INTERCONNECT SplitCLK_4_239_DFFT_84__FPB_n276(net210_c1,net210);
INTERCONNECT SplitCLK_4_238_DFFT_67__FPB_n259(net211_c1,net211);
INTERCONNECT SplitCLK_2_237_DFFT_81__FPB_n273(net212_c1,net212);
INTERCONNECT SplitCLK_4_236_DFFT_63__FPB_n255(net213_c1,net213);
INTERCONNECT SplitCLK_2_235_DFFT_106__FPB_n298(net214_c1,net214);
INTERCONNECT SplitCLK_4_234_DFFT_121__FPB_n313(net215_c1,net215);
INTERCONNECT SplitCLK_2_233_DFFT_112__FPB_n304(net216_c1,net216);
INTERCONNECT SplitCLK_4_232_NOTT_18_n33(net217_c1,net217);
INTERCONNECT SplitCLK_2_231_OR2T_31_n46(net218_c1,net218);
INTERCONNECT SplitCLK_2_230_AND2T_43_n58(net219_c1,net219);
INTERCONNECT SplitCLK_4_229_AND2T_50_n65(net220_c1,net220);
INTERCONNECT SplitCLK_4_228_AND2T_26_n41(net221_c1,net221);
INTERCONNECT SplitCLK_2_227_AND2T_22_n37(net222_c1,net222);
INTERCONNECT SplitCLK_2_226_SplitCLK_6_198(net223_c1,net223);
INTERCONNECT SplitCLK_2_226_SplitCLK_4_225(net224_c1,net224);
INTERCONNECT SplitCLK_4_225_SplitCLK_0_211(net225_c1,net225);
INTERCONNECT SplitCLK_4_225_SplitCLK_2_224(net226_c1,net226);
INTERCONNECT SplitCLK_2_224_SplitCLK_6_217(net227_c1,net227);
INTERCONNECT SplitCLK_2_224_SplitCLK_4_223(net228_c1,net228);
INTERCONNECT SplitCLK_4_223_SplitCLK_4_220(net229_c1,net229);
INTERCONNECT SplitCLK_4_223_SplitCLK_2_222(net230_c1,net230);
INTERCONNECT SplitCLK_2_222_SplitCLK_4_238(net231_c1,net231);
INTERCONNECT SplitCLK_2_222_SplitCLK_4_221(net232_c1,net232);
INTERCONNECT SplitCLK_4_221_OR2T_11_n26(net233_c1,net233);
INTERCONNECT SplitCLK_4_221_DFFT_68__FPB_n260(net234_c1,net234);
INTERCONNECT SplitCLK_4_220_SplitCLK_4_218(net235_c1,net235);
INTERCONNECT SplitCLK_4_220_SplitCLK_4_219(net236_c1,net236);
INTERCONNECT SplitCLK_4_219_AND2T_29_n44(net237_c1,net237);
INTERCONNECT SplitCLK_4_219_DFFT_58__FBL_n250(net238_c1,net238);
INTERCONNECT SplitCLK_4_218_AND2T_17_n32(net239_c1,net239);
INTERCONNECT SplitCLK_4_218_DFFT_79__FPB_n271(net240_c1,net240);
INTERCONNECT SplitCLK_6_217_SplitCLK_0_214(net241_c1,net241);
INTERCONNECT SplitCLK_6_217_SplitCLK_2_216(net242_c1,net242);
INTERCONNECT SplitCLK_2_216_SplitCLK_4_234(net243_c1,net243);
INTERCONNECT SplitCLK_2_216_SplitCLK_4_215(net244_c1,net244);
INTERCONNECT SplitCLK_4_215_AND2T_57_n72(net245_c1,net245);
INTERCONNECT SplitCLK_4_215_OR2T_39_n54(net246_c1,net246);
INTERCONNECT SplitCLK_0_214_SplitCLK_0_212(net247_c1,net247);
INTERCONNECT SplitCLK_0_214_SplitCLK_4_213(net248_c1,net248);
INTERCONNECT SplitCLK_4_213_OR2T_25_n40(net249_c1,net249);
INTERCONNECT SplitCLK_4_213_DFFT_91__FPB_n283(net250_c1,net250);
INTERCONNECT SplitCLK_0_212_AND2T_40_n55(net251_c1,net251);
INTERCONNECT SplitCLK_0_212_DFFT_90__FPB_n282(net252_c1,net252);
INTERCONNECT SplitCLK_0_211_SplitCLK_2_204(net253_c1,net253);
INTERCONNECT SplitCLK_0_211_SplitCLK_4_210(net254_c1,net254);
INTERCONNECT SplitCLK_4_210_SplitCLK_0_207(net255_c1,net255);
INTERCONNECT SplitCLK_4_210_SplitCLK_2_209(net256_c1,net256);
INTERCONNECT SplitCLK_2_209_SplitCLK_4_239(net257_c1,net257);
INTERCONNECT SplitCLK_2_209_SplitCLK_4_208(net258_c1,net258);
INTERCONNECT SplitCLK_4_208_NOTT_9_n24(net259_c1,net259);
INTERCONNECT SplitCLK_4_208_OR2T_28_n43(net260_c1,net260);
INTERCONNECT SplitCLK_0_207_SplitCLK_4_205(net261_c1,net261);
INTERCONNECT SplitCLK_0_207_SplitCLK_4_206(net262_c1,net262);
INTERCONNECT SplitCLK_4_206_DFFT_82__FPB_n274(net263_c1,net263);
INTERCONNECT SplitCLK_4_206_DFFT_83__FPB_n275(net264_c1,net264);
INTERCONNECT SplitCLK_4_205_OR2T_27_n42(net265_c1,net265);
INTERCONNECT SplitCLK_4_205_DFFT_76__FPB_n268(net266_c1,net266);
INTERCONNECT SplitCLK_2_204_SplitCLK_0_201(net267_c1,net267);
INTERCONNECT SplitCLK_2_204_SplitCLK_2_203(net268_c1,net268);
INTERCONNECT SplitCLK_2_203_SplitCLK_4_228(net269_c1,net269);
INTERCONNECT SplitCLK_2_203_SplitCLK_4_202(net270_c1,net270);
INTERCONNECT SplitCLK_4_202_OR2T_33_n48(net271_c1,net271);
INTERCONNECT SplitCLK_4_202_DFFT_78__FPB_n270(net272_c1,net272);
INTERCONNECT SplitCLK_0_201_SplitCLK_4_199(net273_c1,net273);
INTERCONNECT SplitCLK_0_201_SplitCLK_4_200(net274_c1,net274);
INTERCONNECT SplitCLK_4_200_OR2T_34_n49(net275_c1,net275);
INTERCONNECT SplitCLK_4_200_DFFT_75__FPB_n267(net276_c1,net276);
INTERCONNECT SplitCLK_4_199_AND2T_35_n50(net277_c1,net277);
INTERCONNECT SplitCLK_4_199_AND2T_36_n51(net278_c1,net278);
INTERCONNECT SplitCLK_6_198_SplitCLK_0_184(net279_c1,net279);
INTERCONNECT SplitCLK_6_198_SplitCLK_2_197(net280_c1,net280);
INTERCONNECT SplitCLK_2_197_SplitCLK_6_190(net281_c1,net281);
INTERCONNECT SplitCLK_2_197_SplitCLK_4_196(net282_c1,net282);
INTERCONNECT SplitCLK_4_196_SplitCLK_0_193(net283_c1,net283);
INTERCONNECT SplitCLK_4_196_SplitCLK_2_195(net284_c1,net284);
INTERCONNECT SplitCLK_2_195_SplitCLK_2_235(net285_c1,net285);
INTERCONNECT SplitCLK_2_195_SplitCLK_4_194(net286_c1,net286);
INTERCONNECT SplitCLK_4_194_DFFT_99__FPB_n291(net287_c1,net287);
INTERCONNECT SplitCLK_4_194_OR2T_45_n60(net288_c1,net288);
INTERCONNECT SplitCLK_0_193_SplitCLK_0_191(net289_c1,net289);
INTERCONNECT SplitCLK_0_193_SplitCLK_4_192(net290_c1,net290);
INTERCONNECT SplitCLK_4_192_DFFT_111__FPB_n303(net291_c1,net291);
INTERCONNECT SplitCLK_4_192_DFFT_89__FPB_n281(net292_c1,net292);
INTERCONNECT SplitCLK_0_191_AND2T_46_n61(net293_c1,net293);
INTERCONNECT SplitCLK_0_191_OR2T_44_n59(net294_c1,net294);
INTERCONNECT SplitCLK_6_190_SplitCLK_4_187(net295_c1,net295);
INTERCONNECT SplitCLK_6_190_SplitCLK_2_189(net296_c1,net296);
INTERCONNECT SplitCLK_2_189_SplitCLK_4_240(net297_c1,net297);
INTERCONNECT SplitCLK_2_189_SplitCLK_4_188(net298_c1,net298);
INTERCONNECT SplitCLK_4_188_DFFT_65__FPB_n257(net299_c1,net299);
INTERCONNECT SplitCLK_4_188_DFFT_74__FPB_n266(net300_c1,net300);
INTERCONNECT SplitCLK_4_187_SplitCLK_0_185(net301_c1,net301);
INTERCONNECT SplitCLK_4_187_SplitCLK_4_186(net302_c1,net302);
INTERCONNECT SplitCLK_4_186_AND2T_23_n38(net303_c1,net303);
INTERCONNECT SplitCLK_4_186_DFFT_60__FBL_n252(net304_c1,net304);
INTERCONNECT SplitCLK_0_185_DFFT_118__FPB_n310(net305_c1,net305);
INTERCONNECT SplitCLK_0_185_DFFT_62__FBL_n254(net306_c1,net306);
INTERCONNECT SplitCLK_0_184_SplitCLK_6_177(net307_c1,net307);
INTERCONNECT SplitCLK_0_184_SplitCLK_4_183(net308_c1,net308);
INTERCONNECT SplitCLK_4_183_SplitCLK_0_180(net309_c1,net309);
INTERCONNECT SplitCLK_4_183_SplitCLK_2_182(net310_c1,net310);
INTERCONNECT SplitCLK_2_182_SplitCLK_2_230(net311_c1,net311);
INTERCONNECT SplitCLK_2_182_SplitCLK_4_181(net312_c1,net312);
INTERCONNECT SplitCLK_4_181_AND2T_41_n56(net313_c1,net313);
INTERCONNECT SplitCLK_4_181_DFFT_100__FPB_n292(net314_c1,net314);
INTERCONNECT SplitCLK_0_180_SplitCLK_4_178(net315_c1,net315);
INTERCONNECT SplitCLK_0_180_SplitCLK_4_179(net316_c1,net316);
INTERCONNECT SplitCLK_4_179_AND2T_21_n36(net317_c1,net317);
INTERCONNECT SplitCLK_4_179_DFFT_59__FBL_n251(net318_c1,net318);
INTERCONNECT SplitCLK_4_178_OR2T_42_n57(net319_c1,net319);
INTERCONNECT SplitCLK_4_178_DFFT_105__FPB_n297(net320_c1,net320);
INTERCONNECT SplitCLK_6_177_SplitCLK_4_173(net321_c1,net321);
INTERCONNECT SplitCLK_6_177_SplitCLK_6_176(net322_c1,net322);
INTERCONNECT SplitCLK_6_176_SplitCLK_0_174(net323_c1,net323);
INTERCONNECT SplitCLK_6_176_SplitCLK_4_175(net324_c1,net324);
INTERCONNECT SplitCLK_4_175_NOTT_13_n28(net325_c1,net325);
INTERCONNECT SplitCLK_4_175_DFFT_102__FPB_n294(net326_c1,net326);
INTERCONNECT SplitCLK_0_174_NOTT_14_n29(net327_c1,net327);
INTERCONNECT SplitCLK_0_174_DFFT_119__FPB_n311(net328_c1,net328);
INTERCONNECT SplitCLK_4_173_SplitCLK_4_171(net329_c1,net329);
INTERCONNECT SplitCLK_4_173_SplitCLK_4_172(net330_c1,net330);
INTERCONNECT SplitCLK_4_172_AND2T_15_n30(net331_c1,net331);
INTERCONNECT SplitCLK_4_172_DFFT_101__FPB_n293(net332_c1,net332);
INTERCONNECT SplitCLK_4_171_XOR2T_55_n70(net333_c1,net333);
INTERCONNECT SplitCLK_4_171_DFFT_70__FPB_n262(net334_c1,net334);
INTERCONNECT SplitCLK_0_170_SplitCLK_6_142(net335_c1,net335);
INTERCONNECT SplitCLK_0_170_SplitCLK_4_169(net336_c1,net336);
INTERCONNECT SplitCLK_4_169_SplitCLK_0_155(net337_c1,net337);
INTERCONNECT SplitCLK_4_169_SplitCLK_4_168(net338_c1,net338);
INTERCONNECT SplitCLK_4_168_SplitCLK_6_161(net339_c1,net339);
INTERCONNECT SplitCLK_4_168_SplitCLK_4_167(net340_c1,net340);
INTERCONNECT SplitCLK_4_167_SplitCLK_0_164(net341_c1,net341);
INTERCONNECT SplitCLK_4_167_SplitCLK_6_166(net342_c1,net342);
INTERCONNECT SplitCLK_6_166_SplitCLK_2_237(net343_c1,net343);
INTERCONNECT SplitCLK_6_166_SplitCLK_4_165(net344_c1,net344);
INTERCONNECT SplitCLK_4_165_DFFT_80__FPB_n272(net345_c1,net345);
INTERCONNECT SplitCLK_4_165_DFFT_77__FPB_n269(net346_c1,net346);
INTERCONNECT SplitCLK_0_164_SplitCLK_0_162(net347_c1,net347);
INTERCONNECT SplitCLK_0_164_SplitCLK_4_163(net348_c1,net348);
INTERCONNECT SplitCLK_4_163_NOTT_8_n23(net349_c1,net349);
INTERCONNECT SplitCLK_4_163_DFFT_93__FPB_n285(net350_c1,net350);
INTERCONNECT SplitCLK_0_162_DFFT_71__FPB_n263(net351_c1,net351);
INTERCONNECT SplitCLK_0_162_DFFT_72__FPB_n264(net352_c1,net352);
INTERCONNECT SplitCLK_6_161_SplitCLK_0_158(net353_c1,net353);
INTERCONNECT SplitCLK_6_161_SplitCLK_6_160(net354_c1,net354);
INTERCONNECT SplitCLK_6_160_SplitCLK_4_232(net355_c1,net355);
INTERCONNECT SplitCLK_6_160_SplitCLK_4_159(net356_c1,net356);
INTERCONNECT SplitCLK_4_159_AND2T_24_n39(net357_c1,net357);
INTERCONNECT SplitCLK_4_159_OR2T_19_n34(net358_c1,net358);
INTERCONNECT SplitCLK_0_158_SplitCLK_0_156(net359_c1,net359);
INTERCONNECT SplitCLK_0_158_SplitCLK_4_157(net360_c1,net360);
INTERCONNECT SplitCLK_4_157_AND2T_10_n25(net361_c1,net361);
INTERCONNECT SplitCLK_4_157_DFFT_66__FPB_n258(net362_c1,net362);
INTERCONNECT SplitCLK_0_156_AND2T_16_n31(net363_c1,net363);
INTERCONNECT SplitCLK_0_156_DFFT_92__FPB_n284(net364_c1,net364);
INTERCONNECT SplitCLK_0_155_SplitCLK_4_148(net365_c1,net365);
INTERCONNECT SplitCLK_0_155_SplitCLK_4_154(net366_c1,net366);
INTERCONNECT SplitCLK_4_154_SplitCLK_4_151(net367_c1,net367);
INTERCONNECT SplitCLK_4_154_SplitCLK_2_153(net368_c1,net368);
INTERCONNECT SplitCLK_2_153_SplitCLK_2_227(net369_c1,net369);
INTERCONNECT SplitCLK_2_153_SplitCLK_4_152(net370_c1,net370);
INTERCONNECT SplitCLK_4_152_OR2T_12_n27(net371_c1,net371);
INTERCONNECT SplitCLK_4_152_DFFT_73__FPB_n265(net372_c1,net372);
INTERCONNECT SplitCLK_4_151_SplitCLK_4_149(net373_c1,net373);
INTERCONNECT SplitCLK_4_151_SplitCLK_4_150(net374_c1,net374);
INTERCONNECT SplitCLK_4_150_DFFT_94__FPB_n286(net375_c1,net375);
INTERCONNECT SplitCLK_4_150_DFFT_96__FPB_n288(net376_c1,net376);
INTERCONNECT SplitCLK_4_149_DFFT_69__FPB_n261(net377_c1,net377);
INTERCONNECT SplitCLK_4_149_DFFT_95__FPB_n287(net378_c1,net378);
INTERCONNECT SplitCLK_4_148_SplitCLK_6_145(net379_c1,net379);
INTERCONNECT SplitCLK_4_148_SplitCLK_2_147(net380_c1,net380);
INTERCONNECT SplitCLK_2_147_SplitCLK_2_233(net381_c1,net381);
INTERCONNECT SplitCLK_2_147_SplitCLK_4_146(net382_c1,net382);
INTERCONNECT SplitCLK_4_146_AND2T_38_n53(net383_c1,net383);
INTERCONNECT SplitCLK_4_146_DFFT_107__FPB_n299(net384_c1,net384);
INTERCONNECT SplitCLK_6_145_SplitCLK_4_143(net385_c1,net385);
INTERCONNECT SplitCLK_6_145_SplitCLK_4_144(net386_c1,net386);
INTERCONNECT SplitCLK_4_144_DFFT_108__FPB_n300(net387_c1,net387);
INTERCONNECT SplitCLK_4_144_DFFT_97__FPB_n289(net388_c1,net388);
INTERCONNECT SplitCLK_4_143_DFFT_110__FPB_n302(net389_c1,net389);
INTERCONNECT SplitCLK_4_143_DFFT_109__FPB_n301(net390_c1,net390);
INTERCONNECT SplitCLK_6_142_SplitCLK_0_128(net391_c1,net391);
INTERCONNECT SplitCLK_6_142_SplitCLK_6_141(net392_c1,net392);
INTERCONNECT SplitCLK_6_141_SplitCLK_6_134(net393_c1,net393);
INTERCONNECT SplitCLK_6_141_SplitCLK_6_140(net394_c1,net394);
INTERCONNECT SplitCLK_6_140_SplitCLK_0_137(net395_c1,net395);
INTERCONNECT SplitCLK_6_140_SplitCLK_2_139(net396_c1,net396);
INTERCONNECT SplitCLK_2_139_SplitCLK_4_229(net397_c1,net397);
INTERCONNECT SplitCLK_2_139_SplitCLK_4_138(net398_c1,net398);
INTERCONNECT SplitCLK_4_138_AND2T_20_n35(net399_c1,net399);
INTERCONNECT SplitCLK_4_138_DFFT_61__FBL_n253(net400_c1,net400);
INTERCONNECT SplitCLK_0_137_SplitCLK_4_135(net401_c1,net401);
INTERCONNECT SplitCLK_0_137_SplitCLK_4_136(net402_c1,net402);
INTERCONNECT SplitCLK_4_136_AND2T_30_n45(net403_c1,net403);
INTERCONNECT SplitCLK_4_136_OR2T_51_n66(net404_c1,net404);
INTERCONNECT SplitCLK_4_135_DFFT_103__FPB_n295(net405_c1,net405);
INTERCONNECT SplitCLK_4_135_DFFT_104__FPB_n296(net406_c1,net406);
INTERCONNECT SplitCLK_6_134_SplitCLK_0_131(net407_c1,net407);
INTERCONNECT SplitCLK_6_134_SplitCLK_2_133(net408_c1,net408);
INTERCONNECT SplitCLK_2_133_SplitCLK_4_236(net409_c1,net409);
INTERCONNECT SplitCLK_2_133_SplitCLK_4_132(net410_c1,net410);
INTERCONNECT SplitCLK_4_132_AND2T_54_n69(net411_c1,net411);
INTERCONNECT SplitCLK_4_132_DFFT_64__FPB_n256(net412_c1,net412);
INTERCONNECT SplitCLK_0_131_SplitCLK_0_129(net413_c1,net413);
INTERCONNECT SplitCLK_0_131_SplitCLK_4_130(net414_c1,net414);
INTERCONNECT SplitCLK_4_130_AND2T_53_n68(net415_c1,net415);
INTERCONNECT SplitCLK_4_130_OR2T_47_n62(net416_c1,net416);
INTERCONNECT SplitCLK_0_129_AND2T_56_n71(net417_c1,net417);
INTERCONNECT SplitCLK_0_129_DFFT_117__FPB_n309(net418_c1,net418);
INTERCONNECT SplitCLK_0_128_SplitCLK_6_121(net419_c1,net419);
INTERCONNECT SplitCLK_0_128_SplitCLK_4_127(net420_c1,net420);
INTERCONNECT SplitCLK_4_127_SplitCLK_0_124(net421_c1,net421);
INTERCONNECT SplitCLK_4_127_SplitCLK_6_126(net422_c1,net422);
INTERCONNECT SplitCLK_6_126_SplitCLK_2_231(net423_c1,net423);
INTERCONNECT SplitCLK_6_126_SplitCLK_4_125(net424_c1,net424);
INTERCONNECT SplitCLK_4_125_AND2T_49_n64(net425_c1,net425);
INTERCONNECT SplitCLK_4_125_OR2T_37_n52(net426_c1,net426);
INTERCONNECT SplitCLK_0_124_SplitCLK_0_122(net427_c1,net427);
INTERCONNECT SplitCLK_0_124_SplitCLK_4_123(net428_c1,net428);
INTERCONNECT SplitCLK_4_123_AND2T_32_n47(net429_c1,net429);
INTERCONNECT SplitCLK_4_123_DFFT_88__FPB_n280(net430_c1,net430);
INTERCONNECT SplitCLK_0_122_DFFT_86__FPB_n278(net431_c1,net431);
INTERCONNECT SplitCLK_0_122_DFFT_87__FPB_n279(net432_c1,net432);
INTERCONNECT SplitCLK_6_121_SplitCLK_4_117(net433_c1,net433);
INTERCONNECT SplitCLK_6_121_SplitCLK_2_120(net434_c1,net434);
INTERCONNECT SplitCLK_2_120_SplitCLK_4_118(net435_c1,net435);
INTERCONNECT SplitCLK_2_120_SplitCLK_4_119(net436_c1,net436);
INTERCONNECT SplitCLK_4_119_OR2T_52_n67(net437_c1,net437);
INTERCONNECT SplitCLK_4_119_DFFT_113__FPB_n305(net438_c1,net438);
INTERCONNECT SplitCLK_4_118_AND2T_48_n63(net439_c1,net439);
INTERCONNECT SplitCLK_4_118_DFFT_116__FPB_n308(net440_c1,net440);
INTERCONNECT SplitCLK_4_117_SplitCLK_4_115(net441_c1,net441);
INTERCONNECT SplitCLK_4_117_SplitCLK_4_116(net442_c1,net442);
INTERCONNECT SplitCLK_4_116_DFFT_115__FPB_n307(net443_c1,net443);
INTERCONNECT SplitCLK_4_116_DFFT_85__FPB_n277(net444_c1,net444);
INTERCONNECT SplitCLK_4_115_DFFT_120__FPB_n312(net445_c1,net445);
INTERCONNECT SplitCLK_4_115_DFFT_114__FPB_n306(net446_c1,net446);
INTERCONNECT GCLK_Pad_SplitCLK_0_241(GCLK_Pad,net447);
INTERCONNECT Split_HOLD_294_DFFT_101__FPB_n293(net448_c1,net448);
INTERCONNECT Split_HOLD_295_AND2T_26_n41(net449_c1,net449);

endmodule
