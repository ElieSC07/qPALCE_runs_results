// Verilog for Boundary Scan Architecture of Figure 10-15
module TAP(clk, TMS, TDO, St_obs0, St_obs1, St_obs2);

    input clk, TMS;
    output TDO, St_obs0, St_obs1, St_obs2;                     
    reg TDO, St_obs0, St_obs1, St_obs2; 
    reg[3:0] St;

    //TAP Controller States
    parameter[3:0] TestLogicReset = 0, RunTestIdle = 1, SelectDRScan = 2, CaptureDR = 3, ShiftDR = 4, Exit1DR = 5, PauseDR = 6, Exit2DR = 7, UpdateDR = 8, SelectIRScan = 9, CaptureIR = 10, ShiftIR = 11, Exit1IR = 12, PauseIR = 13, Exit2IR = 14, UpdateIR = 15; 
    
    //assign TDO = 0;

    always @(posedge clk)
        begin
            case (St)
                TestLogicReset :
                    begin
                    if (TMS == 1'b0)
                        St <= RunTestIdle ;
                    else
                        St <= TestLogicReset ;
                    end

                RunTestIdle :
                    begin
                        if (TMS == 1'b0)
                            St <= RunTestIdle ;
                        else
                            st <= SelectDRScan ;
                    end

                SelectDRScan :
                    begin 
                        if (TMS == 1'b0)
                            St <= CaptureDR ;
                        else
                            St <= SelectIRScan ;
                    end

                CaptureDR:
                    begin
                        if (TMS == 1'b0)
                            St <= ShiftDR ; 
                        else
                            St <= Exit1DR ;
                    end
    
                ShiftDR:
                    begin
                        if (TMS == 1'b0)
                            St <= ShiftDR ;
                        else
                            St <= Exit1DR ;
                    end

                Exit1DR :
                    begin
                        if (TMS == 1'b0)
                            St <= PauseDR ;
                        else
                            St <= UpdateDR ;
                    end

                PauseDR :
                    begin
                        if (TMS == 1'b0)
                            St <= PauseDR ;
                        else
                            St <= Exit2DR ;
                    end

                Exit2DR :
                    begin
                        if (TMS == 1'b0)
                            St <= ShiftDR ;
                        else
                            st <= UpdateDR ;
                    end

                UpdateDR :
                    begin
                        if (TMS == 1'b0)
                            St <= RunTestIdle ;
                        else
                            St <= SelectDRScan ;
                    end

                SelectIRScan :
                    begin
                        if (TMS == 1'b0)
                            St <= CaptureIR ;
                        else
                            St <= TestLogicReset ;
                    end

                CaptureIR :
                    begin
                        if (TMS == 1'b0)
                            St <= ShiftIR ;
                        else
                            St <= Exit1IR ;
                    end

                ShiftIR: 
                    begin
                        if (TMS == 1'b0)
                            St <= ShiftIR ;
                        else
                            St <= Exit1IR ;
                    end

                Exit1IR :
                    begin
                        if (TMS == 1'b0)
                            St <= PauseIR ;
                        else
                            St <= UpdateIR ;
                    end

                PauseIR :
                    begin
                        if (TMS == 1'b0)
                            St <= PauseIR ;
                        else
                            St <= Exit2IR ;
                    end

                Exit2IR:
                    begin
                        if (TMS == 1'b0)
                            St <= ShiftIR ;
                        else
                            St <= UpdateIR ;
                    end

                UpdateIR:
                    begin
                        if (TMS == 1'b0)
                            St <= RunTestIdle ;
                        else
                            St <= SelectDRScan ;
                    end
            endcase
        end

   always @(St)
    begin
        if ( St == TestLogicReset ) begin
            TDO <= 1'b1;
            St_obs0 <= 1'b1; 
            St_obs1 <= 1'b1;  
            St_obs2 <= 1'b1;
        end
        else begin
            TDO <= 1'b0; 
            St_obs0 <= 1'b0; 
            St_obs1 <= 1'b0;  
            St_obs2 <= 1'b0;
        end
    end

endmodule














