module TAP_half_route(
input GCLK_Pad,
input TMS_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output state_obs2_Pad,
output state_obs3_Pad);

wire TMS_Pad;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire TRST_Pad;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire state_obs0_Pad;
wire net229_c1;
wire state_obs1_Pad;
wire net230_c1;
wire state_obs2_Pad;
wire net231_c1;
wire state_obs3_Pad;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire GCLK_Pad;
wire net486;

DFFT DFFT_99__FPB_n300(net250,net128,net179_c1);
XOR2T XOR2T_29_n65(net344,net160,net153,net24_c1);
DFFT DFFT_63_state_obs0_buf(net326,net169,net161_c1);
DFFT DFFT_64_state_obs1_buf(net350,net170,net162_c1);
DFFT DFFT_65_state_obs2_buf(net448,net171,net163_c1);
DFFT DFFT_66_state_obs3_buf(net478,net172,net164_c1);
AND2T AND2T_9_n45(net314,net145,net217,net8_c1);
NOTT NOTT_8_n44(net476,net142,net5_c1);
AND2T AND2T_10_n46(net338,net94,net219,net12_c1);
AND2T AND2T_11_n47(net336,net149,net221,net16_c1);
AND2T AND2T_20_n56(net308,net98,net75,net20_c1);
AND2T AND2T_21_n57(net432,net115,net225,net25_c1);
AND2T AND2T_14_n50(net462,net117,net113,net1_c1);
AND2T AND2T_30_n66(net440,net66,net216,net30_c1);
AND2T AND2T_22_n58(net470,net70,net132,net31_c1);
AND2T AND2T_31_n67(net434,net30,net112,net35_c1);
AND2T AND2T_24_n60(net468,net80,net212,net3_c1);
AND2T AND2T_16_n52(net315,net125,net223,net4_c1);
AND2T AND2T_40_n76(net372,net34,net110,net39_c1);
AND2T AND2T_25_n61(net296,net63,net213,net6_c1);
AND2T AND2T_17_n53(net345,net4,net120,net7_c1);
AND2T AND2T_50_n86(net276,net78,net187,net46_c1);
AND2T AND2T_35_n71(net414,net116,net227,net13_c1);
AND2T AND2T_19_n55(net312,net106,net97,net15_c1);
AND2T AND2T_51_n87(net264,net46,net38,net49_c1);
AND2T AND2T_43_n79(net258,net47,net23,net50_c1);
AND2T AND2T_44_n80(net260,net127,net194,net17_c1);
AND2T AND2T_28_n64(net446,net137,net215,net19_c1);
AND2T AND2T_60_n96(net384,net48,net58,net51_c1);
AND2T AND2T_45_n81(net288,net93,net198,net22_c1);
AND2T AND2T_61_n97(net385,net51,net207,net53_c1);
AND2T AND2T_53_n89(net259,net52,net72,net54_c1);
AND2T AND2T_54_n90(net420,net74,net197,net27_c1);
AND2T AND2T_46_n82(net378,net140,net202,net28_c1);
AND2T AND2T_62_n98(net416,net65,net186,net55_c1);
AND2T AND2T_47_n83(net390,net130,net204,net33_c1);
AND2T AND2T_39_n75(net282,net61,net184,net34_c1);
AND2T AND2T_57_n93(net417,net122,net201,net41_c1);
AND2T AND2T_59_n95(net280,net134,net203,net48_c1);
OR2T OR2T_23_n59(net438,net31,net25,net36_c1);
OR2T OR2T_32_n68(net433,net35,net129,net40_c1);
OR2T OR2T_41_n77(net391,net39,net190,net43_c1);
OR2T OR2T_33_n69(net266,net147,net218,net44_c1);
OR2T OR2T_34_n70(net392,net44,net14,net9_c1);
OR2T OR2T_26_n62(net408,net135,net126,net10_c1);
OR2T OR2T_42_n78(net294,net144,net69,net47_c1);
OR2T OR2T_27_n63(net393,net10,net121,net14_c1);
OR2T OR2T_36_n72(net370,net85,net182,net18_c1);
OR2T OR2T_52_n88(net246,net49,net189,net52_c1);
OR2T OR2T_37_n73(net277,net131,net96,net23_c1);
OR2T OR2T_55_n91(net415,net27,net118,net32_c1);
OR2T OR2T_56_n92(net421,net32,net151,net37_c1);
OR2T OR2T_48_n84(net295,net33,net143,net38_c1);
OR2T OR2T_49_n85(net244,net155,net73,net42_c1);
NOTT NOTT_12_n48(net313,net150,net21_c1);
NOTT NOTT_13_n49(net342,net158,net26_c1);
NOTT NOTT_15_n51(net435,net159,net2_c1);
NOTT NOTT_18_n54(net402,net107,net11_c1);
NOTT NOTT_38_n74(net281,net124,net29_c1);
NOTT NOTT_58_n94(net290,net114,net45_c1);
AND2T AND2T_67_n109(net477,net5,net188,net57_c1);
DFFT DFFT_100__FPB_n301(net274,net179,net180_c1);
DFFT DFFT_101__FPB_n302(net275,net180,net182_c1);
DFFT DFFT_110__FPB_n311(net252,net181,net183_c1);
DFFT DFFT_102__FPB_n303(net283,net104,net184_c1);
DFFT DFFT_111__FPB_n312(net253,net183,net187_c1);
DFFT DFFT_103__FPB_n304(net403,net89,net185_c1);
DFFT DFFT_70__PIPL_n112(net356,net162,net166_c1);
DFFT DFFT_120__FPB_n321(net464,net157,net188_c1);
DFFT DFFT_112__FPB_n313(net265,net100,net189_c1);
DFFT DFFT_104__FPB_n305(net409,net185,net190_c1);
DFFT DFFT_121__FPB_n322(net320,net165,net192_c1);
DFFT DFFT_113__FPB_n314(net406,net136,net193_c1);
DFFT DFFT_105__FPB_n306(net261,net50,net194_c1);
DFFT DFFT_71__PIPL_n113(net452,net163,net167_c1);
DFFT DFFT_130__FPB_n331(net449,net191,net195_c1);
DFFT DFFT_122__FPB_n323(net328,net192,net196_c1);
DFFT DFFT_114__FPB_n315(net407,net193,net197_c1);
DFFT DFFT_106__FPB_n307(net291,net87,net198_c1);
DFFT DFFT_131__FPB_n332(net358,net195,net199_c1);
DFFT DFFT_123__FPB_n324(net322,net196,net200_c1);
DFFT DFFT_115__FPB_n316(net422,net37,net201_c1);
DFFT DFFT_107__FPB_n308(net373,net152,net202_c1);
DFFT DFFT_72__PIPL_n114(net482,net164,net168_c1);
DFFT DFFT_116__FPB_n317(net251,net76,net203_c1);
DFFT DFFT_108__FPB_n309(net379,net28,net204_c1);
DFFT DFFT_109__FPB_n310(net245,net42,net181_c1);
DFFT DFFT_133__FPB_n334(net484,net168,net205_c1);
DFFT DFFT_125__FPB_n326(net357,net166,net206_c1);
DFFT DFFT_117__FPB_n318(net297,net45,net207_c1);
DFFT DFFT_73__PIPL_n115(net327,net8,net169_c1);
DFFT DFFT_134__FPB_n335(net485,net205,net208_c1);
DFFT DFFT_126__FPB_n327(net352,net206,net209_c1);
DFFT DFFT_118__FPB_n319(net386,net53,net210_c1);
DFFT DFFT_119__FPB_n320(net387,net210,net186_c1);
DFFT DFFT_127__FPB_n328(net353,net209,net211_c1);
DFFT DFFT_74__PIPL_n116(net351,net12,net170_c1);
DFFT DFFT_129__FPB_n330(net454,net167,net191_c1);
DFFT DFFT_75__PIPL_n117(net453,net84,net171_c1);
DFFT DFFT_80__FBL_n281(net471,net214,net174_c1);
DFFT DFFT_76__PIPL_n118(net479,net79,net172_c1);
DFFT DFFT_81__FBL_n282(net306,net95,net175_c1);
DFFT DFFT_124_state_obs0(net323,net200,net228_c1);
DFFT DFFT_132_state_obs2(net359,net199,net230_c1);
DFFT DFFT_82__FBL_n283(net307,net103,net176_c1);
DFFT DFFT_69__PIPL_n111(net321,net161,net165_c1);
DFFT DFFT_90__FPB_n291(net267,net62,net213_c1);
SPLITT Split_140_n341(net21,net59_c1,net111_c1);
SPLITT Split_141_n342(net111,net61_c1,net113_c1);
SPLITT Split_142_n343(net59,net62_c1,net114_c1);
SPLITT Split_150_n351(net60,net63_c1,net115_c1);
SPLITT Split_143_n344(net26,net66_c1,net117_c1);
SPLITT Split_151_n352(net36,net64_c1,net118_c1);
SPLITT Split_136_n337(net0,net67_c1,net119_c1);
SPLITT Split_144_n345(net1,net70_c1,net120_c1);
SPLITT Split_152_n353(net64,net69_c1,net121_c1);
SPLITT Split_160_n361(net13,net68_c1,net122_c1);
SPLITT Split_137_n338(net119,net73_c1,net124_c1);
SPLITT Split_145_n346(net2,net75_c1,net125_c1);
SPLITT Split_153_n354(net3,net74_c1,net126_c1);
SPLITT Split_161_n362(net68,net72_c1,net127_c1);
SPLITT Split_138_n339(net67,net76_c1,net128_c1);
SPLITT Split_146_n347(net7,net79_c1,net129_c1);
SPLITT Split_154_n355(net6,net77_c1,net130_c1);
SPLITT Split_162_n363(net18,net78_c1,net131_c1);
SPLITT Split_170_n371(net123,net80_c1,net132_c1);
SPLITT Split_139_n340(net16,net58_c1,net110_c1);
SPLITT Split_147_n348(net11,net83_c1,net134_c1);
SPLITT Split_155_n356(net77,net85_c1,net135_c1);
SPLITT Split_163_n364(net29,net81_c1,net136_c1);
SPLITT Split_171_n372(net71,net84_c1,net137_c1);
SPLITT Split_148_n349(net15,net88_c1,net138_c1);
SPLITT Split_156_n357(net19,net87_c1,net139_c1);
SPLITT Split_164_n365(net81,net89_c1,net140_c1);
SPLITT Split_172_n373(net56,net86_c1,net141_c1);
SPLITT Split_180_n381(net82,net90_c1,net142_c1);
SPLITT Split_149_n350(net20,net60_c1,net112_c1);
SPLITT Split_157_n358(net40,net92_c1,net143_c1);
SPLITT Split_165_n366(net43,net93_c1,net144_c1);
SPLITT Split_173_n374(net141,net94_c1,net145_c1);
SPLITT Split_181_n382(net175,net91_c1,net146_c1);
SPLITT Split_158_n359(net92,net96_c1,net147_c1);
SPLITT Split_166_n367(net17,net95_c1,net148_c1);
SPLITT Split_174_n375(net86,net98_c1,net149_c1);
SPLITT Split_182_n383(net146,net97_c1,net150_c1);
SPLITT Split_159_n360(net9,net65_c1,net116_c1);
SPLITT Split_167_n368(net22,net100_c1,net151_c1);
SPLITT Split_175_n376(net178,net99_c1,net152_c1);
SPLITT Split_183_n384(net91,net101_c1,net153_c1);
SPLITT Split_168_n369(net54,net103_c1,net154_c1);
SPLITT Split_176_n377(net99,net104_c1,net155_c1);
SPLITT Split_184_n385(net176,net102_c1,net156_c1);
SPLITT Split_169_n370(net57,net71_c1,net123_c1);
SPLITT Split_177_n378(net173,net105_c1,net157_c1);
SPLITT Split_185_n386(net156,net106_c1,net158_c1);
DFFT DFFT_91__FPB_n292(net447,net24,net215_c1);
DFFT DFFT_83__FPB_n284(net469,net55,net214_c1);
SPLITT Split_178_n379(net105,net109_c1,net159_c1);
SPLITT Split_186_n387(net102,net108_c1,net160_c1);
SPLITT Split_179_n380(net174,net82_c1,net133_c1);
DFFT DFFT_92__FPB_n293(net343,net177,net216_c1);
DFFT DFFT_84__FPB_n285(net309,net101,net217_c1);
DFFT DFFT_77__FBL_n278(net337,net148,net177_c1);
DFFT DFFT_93__FPB_n294(net289,net139,net218_c1);
DFFT DFFT_85__FPB_n286(net339,net108,net219_c1);
DFFT DFFT_78__FBL_n279(net247,net154,net178_c1);
DFFT DFFT_94__FPB_n295(net400,net83,net220_c1);
DFFT DFFT_86__FPB_n287(net441,net109,net221_c1);
DFFT DFFT_79__FBL_n280(net423,net41,net173_c1);
DFFT DFFT_95__FPB_n296(net401,net220,net222_c1);
DFFT DFFT_87__FPB_n288(net465,net133,net223_c1);
DFFT DFFT_135_state_obs3(net455,net208,net231_c1);
NOTT NOTT_68_n110(net483,net90,net56_c1);
DFFT DFFT_96__FPB_n297(net371,net222,net224_c1);
DFFT DFFT_88__FPB_n289(net439,net138,net225_c1);
DFFT DFFT_89__FPB_n290(net463,net88,net212_c1);
DFFT DFFT_97__FPB_n298(net376,net224,net226_c1);
DFFT DFFT_128_state_obs1(net329,net211,net229_c1);
DFFT DFFT_98__FPB_n299(net377,net226,net227_c1);
SPLITT SplitCLK_4_129(net480,net484_c1,net485_c1);
SPLITT SplitCLK_4_130(net481,net482_c1,net483_c1);
SPLITT SplitCLK_4_131(net472,net481_c1,net480_c1);
SPLITT SplitCLK_4_132(net474,net479_c1,net478_c1);
SPLITT SplitCLK_4_133(net475,net477_c1,net476_c1);
SPLITT SplitCLK_2_134(net473,net475_c1,net474_c1);
SPLITT SplitCLK_6_135(net456,net472_c1,net473_c1);
SPLITT SplitCLK_4_136(net466,net470_c1,net471_c1);
SPLITT SplitCLK_4_137(net467,net468_c1,net469_c1);
SPLITT SplitCLK_0_138(net458,net466_c1,net467_c1);
SPLITT SplitCLK_0_139(net460,net464_c1,net465_c1);
SPLITT SplitCLK_4_140(net461,net462_c1,net463_c1);
SPLITT SplitCLK_2_141(net459,net461_c1,net460_c1);
SPLITT SplitCLK_4_142(net457,net459_c1,net458_c1);
SPLITT SplitCLK_0_143(net424,net456_c1,net457_c1);
SPLITT SplitCLK_4_144(net450,net455_c1,net454_c1);
SPLITT SplitCLK_4_145(net451,net453_c1,net452_c1);
SPLITT SplitCLK_2_146(net442,net450_c1,net451_c1);
SPLITT SplitCLK_4_147(net444,net448_c1,net449_c1);
SPLITT SplitCLK_4_148(net445,net447_c1,net446_c1);
SPLITT SplitCLK_2_149(net443,net445_c1,net444_c1);
SPLITT SplitCLK_6_150(net426,net442_c1,net443_c1);
SPLITT SplitCLK_4_151(net436,net441_c1,net440_c1);
SPLITT SplitCLK_4_152(net437,net439_c1,net438_c1);
SPLITT SplitCLK_4_153(net428,net436_c1,net437_c1);
SPLITT SplitCLK_4_154(net430,net435_c1,net434_c1);
SPLITT SplitCLK_4_155(net431,net433_c1,net432_c1);
SPLITT SplitCLK_6_156(net429,net431_c1,net430_c1);
SPLITT SplitCLK_4_157(net427,net429_c1,net428_c1);
SPLITT SplitCLK_2_158(net425,net427_c1,net426_c1);
SPLITT SplitCLK_6_159(net360,net424_c1,net425_c1);
SPLITT SplitCLK_0_160(net418,net423_c1,net422_c1);
SPLITT SplitCLK_4_161(net419,net421_c1,net420_c1);
SPLITT SplitCLK_0_162(net410,net418_c1,net419_c1);
SPLITT SplitCLK_0_163(net412,net416_c1,net417_c1);
SPLITT SplitCLK_4_164(net413,net414_c1,net415_c1);
SPLITT SplitCLK_6_165(net411,net413_c1,net412_c1);
SPLITT SplitCLK_4_166(net394,net411_c1,net410_c1);
SPLITT SplitCLK_0_167(net404,net408_c1,net409_c1);
SPLITT SplitCLK_4_168(net405,net406_c1,net407_c1);
SPLITT SplitCLK_0_169(net396,net404_c1,net405_c1);
SPLITT SplitCLK_4_170(net398,net402_c1,net403_c1);
SPLITT SplitCLK_4_171(net399,net401_c1,net400_c1);
SPLITT SplitCLK_4_172(net397,net399_c1,net398_c1);
SPLITT SplitCLK_4_173(net395,net397_c1,net396_c1);
SPLITT SplitCLK_0_174(net362,net394_c1,net395_c1);
SPLITT SplitCLK_0_175(net388,net392_c1,net393_c1);
SPLITT SplitCLK_4_176(net389,net391_c1,net390_c1);
SPLITT SplitCLK_4_177(net380,net388_c1,net389_c1);
SPLITT SplitCLK_0_178(net382,net386_c1,net387_c1);
SPLITT SplitCLK_4_179(net383,net384_c1,net385_c1);
SPLITT SplitCLK_6_180(net381,net382_c1,net383_c1);
SPLITT SplitCLK_2_181(net364,net380_c1,net381_c1);
SPLITT SplitCLK_4_182(net374,net379_c1,net378_c1);
SPLITT SplitCLK_4_183(net375,net376_c1,net377_c1);
SPLITT SplitCLK_0_184(net366,net374_c1,net375_c1);
SPLITT SplitCLK_4_185(net368,net373_c1,net372_c1);
SPLITT SplitCLK_4_186(net369,net370_c1,net371_c1);
SPLITT SplitCLK_6_187(net367,net368_c1,net369_c1);
SPLITT SplitCLK_4_188(net365,net367_c1,net366_c1);
SPLITT SplitCLK_4_189(net363,net364_c1,net365_c1);
SPLITT SplitCLK_4_190(net361,net363_c1,net362_c1);
SPLITT SplitCLK_0_191(net232,net360_c1,net361_c1);
SPLITT SplitCLK_0_192(net354,net358_c1,net359_c1);
SPLITT SplitCLK_4_193(net355,net356_c1,net357_c1);
SPLITT SplitCLK_4_194(net346,net354_c1,net355_c1);
SPLITT SplitCLK_0_195(net348,net352_c1,net353_c1);
SPLITT SplitCLK_4_196(net349,net351_c1,net350_c1);
SPLITT SplitCLK_6_197(net347,net348_c1,net349_c1);
SPLITT SplitCLK_6_198(net330,net346_c1,net347_c1);
SPLITT SplitCLK_4_199(net340,net345_c1,net344_c1);
SPLITT SplitCLK_4_200(net341,net342_c1,net343_c1);
SPLITT SplitCLK_4_201(net332,net340_c1,net341_c1);
SPLITT SplitCLK_0_202(net334,net338_c1,net339_c1);
SPLITT SplitCLK_4_203(net335,net337_c1,net336_c1);
SPLITT SplitCLK_6_204(net333,net335_c1,net334_c1);
SPLITT SplitCLK_4_205(net331,net333_c1,net332_c1);
SPLITT SplitCLK_6_206(net298,net331_c1,net330_c1);
SPLITT SplitCLK_0_207(net324,net328_c1,net329_c1);
SPLITT SplitCLK_4_208(net325,net326_c1,net327_c1);
SPLITT SplitCLK_4_209(net316,net324_c1,net325_c1);
SPLITT SplitCLK_0_210(net318,net322_c1,net323_c1);
SPLITT SplitCLK_4_211(net319,net320_c1,net321_c1);
SPLITT SplitCLK_6_212(net317,net318_c1,net319_c1);
SPLITT SplitCLK_6_213(net300,net316_c1,net317_c1);
SPLITT SplitCLK_4_214(net310,net314_c1,net315_c1);
SPLITT SplitCLK_4_215(net311,net313_c1,net312_c1);
SPLITT SplitCLK_0_216(net302,net310_c1,net311_c1);
SPLITT SplitCLK_4_217(net304,net309_c1,net308_c1);
SPLITT SplitCLK_4_218(net305,net306_c1,net307_c1);
SPLITT SplitCLK_2_219(net303,net305_c1,net304_c1);
SPLITT SplitCLK_6_220(net301,net302_c1,net303_c1);
SPLITT SplitCLK_6_221(net299,net300_c1,net301_c1);
SPLITT SplitCLK_6_222(net234,net298_c1,net299_c1);
SPLITT SplitCLK_0_223(net292,net296_c1,net297_c1);
SPLITT SplitCLK_4_224(net293,net294_c1,net295_c1);
SPLITT SplitCLK_0_225(net284,net292_c1,net293_c1);
SPLITT SplitCLK_4_226(net286,net290_c1,net291_c1);
SPLITT SplitCLK_4_227(net287,net289_c1,net288_c1);
SPLITT SplitCLK_6_228(net285,net286_c1,net287_c1);
SPLITT SplitCLK_6_229(net268,net284_c1,net285_c1);
SPLITT SplitCLK_4_230(net278,net282_c1,net283_c1);
SPLITT SplitCLK_4_231(net279,net281_c1,net280_c1);
SPLITT SplitCLK_4_232(net270,net278_c1,net279_c1);
SPLITT SplitCLK_4_233(net272,net276_c1,net277_c1);
SPLITT SplitCLK_4_234(net273,net274_c1,net275_c1);
SPLITT SplitCLK_2_235(net271,net273_c1,net272_c1);
SPLITT SplitCLK_4_236(net269,net271_c1,net270_c1);
SPLITT SplitCLK_4_237(net236,net269_c1,net268_c1);
SPLITT SplitCLK_4_238(net262,net266_c1,net267_c1);
SPLITT SplitCLK_4_239(net263,net265_c1,net264_c1);
SPLITT SplitCLK_0_240(net254,net262_c1,net263_c1);
SPLITT SplitCLK_4_241(net256,net260_c1,net261_c1);
SPLITT SplitCLK_4_242(net257,net259_c1,net258_c1);
SPLITT SplitCLK_2_243(net255,net257_c1,net256_c1);
SPLITT SplitCLK_6_244(net238,net254_c1,net255_c1);
SPLITT SplitCLK_0_245(net248,net252_c1,net253_c1);
SPLITT SplitCLK_4_246(net249,net251_c1,net250_c1);
SPLITT SplitCLK_0_247(net240,net248_c1,net249_c1);
SPLITT SplitCLK_0_248(net242,net246_c1,net247_c1);
SPLITT SplitCLK_4_249(net243,net244_c1,net245_c1);
SPLITT SplitCLK_6_250(net241,net243_c1,net242_c1);
SPLITT SplitCLK_4_251(net239,net241_c1,net240_c1);
SPLITT SplitCLK_2_252(net237,net239_c1,net238_c1);
SPLITT SplitCLK_4_253(net235,net237_c1,net236_c1);
SPLITT SplitCLK_2_254(net233,net235_c1,net234_c1);
SPLITT SplitCLK_0_255(net486,net232_c1,net233_c1);
INTERCONNECT TMS_Pad_Split_136_n337(TMS_Pad,net0);
INTERCONNECT AND2T_14_n50_Split_144_n345(net1_c1,net1);
INTERCONNECT NOTT_15_n51_Split_145_n346(net2_c1,net2);
INTERCONNECT AND2T_24_n60_Split_153_n354(net3_c1,net3);
INTERCONNECT AND2T_16_n52_AND2T_17_n53(net4_c1,net4);
INTERCONNECT NOTT_8_n44_AND2T_67_n109(net5_c1,net5);
INTERCONNECT AND2T_25_n61_Split_154_n355(net6_c1,net6);
INTERCONNECT AND2T_17_n53_Split_146_n347(net7_c1,net7);
INTERCONNECT AND2T_9_n45_DFFT_73__PIPL_n115(net8_c1,net8);
INTERCONNECT OR2T_34_n70_Split_159_n360(net9_c1,net9);
INTERCONNECT OR2T_26_n62_OR2T_27_n63(net10_c1,net10);
INTERCONNECT NOTT_18_n54_Split_147_n348(net11_c1,net11);
INTERCONNECT AND2T_10_n46_DFFT_74__PIPL_n116(net12_c1,net12);
INTERCONNECT AND2T_35_n71_Split_160_n361(net13_c1,net13);
INTERCONNECT OR2T_27_n63_OR2T_34_n70(net14_c1,net14);
INTERCONNECT AND2T_19_n55_Split_148_n349(net15_c1,net15);
INTERCONNECT AND2T_11_n47_Split_139_n340(net16_c1,net16);
INTERCONNECT AND2T_44_n80_Split_166_n367(net17_c1,net17);
INTERCONNECT OR2T_36_n72_Split_162_n363(net18_c1,net18);
INTERCONNECT AND2T_28_n64_Split_156_n357(net19_c1,net19);
INTERCONNECT AND2T_20_n56_Split_149_n350(net20_c1,net20);
INTERCONNECT NOTT_12_n48_Split_140_n341(net21_c1,net21);
INTERCONNECT AND2T_45_n81_Split_167_n368(net22_c1,net22);
INTERCONNECT OR2T_37_n73_AND2T_43_n79(net23_c1,net23);
INTERCONNECT XOR2T_29_n65_DFFT_91__FPB_n292(net24_c1,net24);
INTERCONNECT AND2T_21_n57_OR2T_23_n59(net25_c1,net25);
INTERCONNECT NOTT_13_n49_Split_143_n344(net26_c1,net26);
INTERCONNECT AND2T_54_n90_OR2T_55_n91(net27_c1,net27);
INTERCONNECT AND2T_46_n82_DFFT_108__FPB_n309(net28_c1,net28);
INTERCONNECT NOTT_38_n74_Split_163_n364(net29_c1,net29);
INTERCONNECT AND2T_30_n66_AND2T_31_n67(net30_c1,net30);
INTERCONNECT AND2T_22_n58_OR2T_23_n59(net31_c1,net31);
INTERCONNECT OR2T_55_n91_OR2T_56_n92(net32_c1,net32);
INTERCONNECT AND2T_47_n83_OR2T_48_n84(net33_c1,net33);
INTERCONNECT AND2T_39_n75_AND2T_40_n76(net34_c1,net34);
INTERCONNECT AND2T_31_n67_OR2T_32_n68(net35_c1,net35);
INTERCONNECT OR2T_23_n59_Split_151_n352(net36_c1,net36);
INTERCONNECT OR2T_56_n92_DFFT_115__FPB_n316(net37_c1,net37);
INTERCONNECT OR2T_48_n84_AND2T_51_n87(net38_c1,net38);
INTERCONNECT AND2T_40_n76_OR2T_41_n77(net39_c1,net39);
INTERCONNECT OR2T_32_n68_Split_157_n358(net40_c1,net40);
INTERCONNECT AND2T_57_n93_DFFT_79__FBL_n280(net41_c1,net41);
INTERCONNECT OR2T_49_n85_DFFT_109__FPB_n310(net42_c1,net42);
INTERCONNECT OR2T_41_n77_Split_165_n366(net43_c1,net43);
INTERCONNECT OR2T_33_n69_OR2T_34_n70(net44_c1,net44);
INTERCONNECT NOTT_58_n94_DFFT_117__FPB_n318(net45_c1,net45);
INTERCONNECT AND2T_50_n86_AND2T_51_n87(net46_c1,net46);
INTERCONNECT OR2T_42_n78_AND2T_43_n79(net47_c1,net47);
INTERCONNECT AND2T_59_n95_AND2T_60_n96(net48_c1,net48);
INTERCONNECT AND2T_51_n87_OR2T_52_n88(net49_c1,net49);
INTERCONNECT AND2T_43_n79_DFFT_105__FPB_n306(net50_c1,net50);
INTERCONNECT AND2T_60_n96_AND2T_61_n97(net51_c1,net51);
INTERCONNECT OR2T_52_n88_AND2T_53_n89(net52_c1,net52);
INTERCONNECT AND2T_61_n97_DFFT_118__FPB_n319(net53_c1,net53);
INTERCONNECT AND2T_53_n89_Split_168_n369(net54_c1,net54);
INTERCONNECT AND2T_62_n98_DFFT_83__FPB_n284(net55_c1,net55);
INTERCONNECT NOTT_68_n110_Split_172_n373(net56_c1,net56);
INTERCONNECT AND2T_67_n109_Split_169_n370(net57_c1,net57);
INTERCONNECT Split_139_n340_AND2T_60_n96(net58_c1,net58);
INTERCONNECT Split_140_n341_Split_142_n343(net59_c1,net59);
INTERCONNECT Split_149_n350_Split_150_n351(net60_c1,net60);
INTERCONNECT Split_141_n342_AND2T_39_n75(net61_c1,net61);
INTERCONNECT Split_142_n343_DFFT_90__FPB_n291(net62_c1,net62);
INTERCONNECT Split_150_n351_AND2T_25_n61(net63_c1,net63);
INTERCONNECT Split_151_n352_Split_152_n353(net64_c1,net64);
INTERCONNECT Split_159_n360_AND2T_62_n98(net65_c1,net65);
INTERCONNECT Split_143_n344_AND2T_30_n66(net66_c1,net66);
INTERCONNECT Split_136_n337_Split_138_n339(net67_c1,net67);
INTERCONNECT Split_160_n361_Split_161_n362(net68_c1,net68);
INTERCONNECT Split_152_n353_OR2T_42_n78(net69_c1,net69);
INTERCONNECT Split_144_n345_AND2T_22_n58(net70_c1,net70);
INTERCONNECT Split_169_n370_Split_171_n372(net71_c1,net71);
INTERCONNECT Split_161_n362_AND2T_53_n89(net72_c1,net72);
INTERCONNECT Split_137_n338_OR2T_49_n85(net73_c1,net73);
INTERCONNECT Split_153_n354_AND2T_54_n90(net74_c1,net74);
INTERCONNECT Split_145_n346_AND2T_20_n56(net75_c1,net75);
INTERCONNECT Split_138_n339_DFFT_116__FPB_n317(net76_c1,net76);
INTERCONNECT Split_154_n355_Split_155_n356(net77_c1,net77);
INTERCONNECT Split_162_n363_AND2T_50_n86(net78_c1,net78);
INTERCONNECT Split_146_n347_DFFT_76__PIPL_n118(net79_c1,net79);
INTERCONNECT Split_170_n371_AND2T_24_n60(net80_c1,net80);
INTERCONNECT Split_163_n364_Split_164_n365(net81_c1,net81);
INTERCONNECT Split_179_n380_Split_180_n381(net82_c1,net82);
INTERCONNECT Split_147_n348_DFFT_94__FPB_n295(net83_c1,net83);
INTERCONNECT Split_171_n372_DFFT_75__PIPL_n117(net84_c1,net84);
INTERCONNECT Split_155_n356_OR2T_36_n72(net85_c1,net85);
INTERCONNECT Split_172_n373_Split_174_n375(net86_c1,net86);
INTERCONNECT Split_156_n357_DFFT_106__FPB_n307(net87_c1,net87);
INTERCONNECT Split_148_n349_DFFT_89__FPB_n290(net88_c1,net88);
INTERCONNECT Split_164_n365_DFFT_103__FPB_n304(net89_c1,net89);
INTERCONNECT Split_180_n381_NOTT_68_n110(net90_c1,net90);
INTERCONNECT Split_181_n382_Split_183_n384(net91_c1,net91);
INTERCONNECT Split_157_n358_Split_158_n359(net92_c1,net92);
INTERCONNECT Split_165_n366_AND2T_45_n81(net93_c1,net93);
INTERCONNECT Split_173_n374_AND2T_10_n46(net94_c1,net94);
INTERCONNECT Split_166_n367_DFFT_81__FBL_n282(net95_c1,net95);
INTERCONNECT Split_158_n359_OR2T_37_n73(net96_c1,net96);
INTERCONNECT Split_182_n383_AND2T_19_n55(net97_c1,net97);
INTERCONNECT Split_174_n375_AND2T_20_n56(net98_c1,net98);
INTERCONNECT Split_175_n376_Split_176_n377(net99_c1,net99);
INTERCONNECT Split_167_n368_DFFT_112__FPB_n313(net100_c1,net100);
INTERCONNECT Split_183_n384_DFFT_84__FPB_n285(net101_c1,net101);
INTERCONNECT Split_184_n385_Split_186_n387(net102_c1,net102);
INTERCONNECT Split_168_n369_DFFT_82__FBL_n283(net103_c1,net103);
INTERCONNECT Split_176_n377_DFFT_102__FPB_n303(net104_c1,net104);
INTERCONNECT Split_177_n378_Split_178_n379(net105_c1,net105);
INTERCONNECT Split_185_n386_AND2T_19_n55(net106_c1,net106);
INTERCONNECT TRST_Pad_NOTT_18_n54(TRST_Pad,net107);
INTERCONNECT Split_186_n387_DFFT_85__FPB_n286(net108_c1,net108);
INTERCONNECT Split_178_n379_DFFT_86__FPB_n287(net109_c1,net109);
INTERCONNECT Split_139_n340_AND2T_40_n76(net110_c1,net110);
INTERCONNECT Split_140_n341_Split_141_n342(net111_c1,net111);
INTERCONNECT Split_149_n350_AND2T_31_n67(net112_c1,net112);
INTERCONNECT Split_141_n342_AND2T_14_n50(net113_c1,net113);
INTERCONNECT Split_142_n343_NOTT_58_n94(net114_c1,net114);
INTERCONNECT Split_150_n351_AND2T_21_n57(net115_c1,net115);
INTERCONNECT Split_159_n360_AND2T_35_n71(net116_c1,net116);
INTERCONNECT Split_143_n344_AND2T_14_n50(net117_c1,net117);
INTERCONNECT Split_151_n352_OR2T_55_n91(net118_c1,net118);
INTERCONNECT Split_136_n337_Split_137_n338(net119_c1,net119);
INTERCONNECT Split_144_n345_AND2T_17_n53(net120_c1,net120);
INTERCONNECT Split_152_n353_OR2T_27_n63(net121_c1,net121);
INTERCONNECT Split_160_n361_AND2T_57_n93(net122_c1,net122);
INTERCONNECT Split_169_n370_Split_170_n371(net123_c1,net123);
INTERCONNECT Split_137_n338_NOTT_38_n74(net124_c1,net124);
INTERCONNECT Split_145_n346_AND2T_16_n52(net125_c1,net125);
INTERCONNECT Split_153_n354_OR2T_26_n62(net126_c1,net126);
INTERCONNECT Split_161_n362_AND2T_44_n80(net127_c1,net127);
INTERCONNECT Split_138_n339_DFFT_99__FPB_n300(net128_c1,net128);
INTERCONNECT Split_146_n347_OR2T_32_n68(net129_c1,net129);
INTERCONNECT Split_154_n355_AND2T_47_n83(net130_c1,net130);
INTERCONNECT Split_162_n363_OR2T_37_n73(net131_c1,net131);
INTERCONNECT Split_170_n371_AND2T_22_n58(net132_c1,net132);
INTERCONNECT Split_179_n380_DFFT_87__FPB_n288(net133_c1,net133);
INTERCONNECT Split_147_n348_AND2T_59_n95(net134_c1,net134);
INTERCONNECT Split_155_n356_OR2T_26_n62(net135_c1,net135);
INTERCONNECT Split_163_n364_DFFT_113__FPB_n314(net136_c1,net136);
INTERCONNECT Split_171_n372_AND2T_28_n64(net137_c1,net137);
INTERCONNECT Split_148_n349_DFFT_88__FPB_n289(net138_c1,net138);
INTERCONNECT Split_156_n357_DFFT_93__FPB_n294(net139_c1,net139);
INTERCONNECT Split_164_n365_AND2T_46_n82(net140_c1,net140);
INTERCONNECT Split_172_n373_Split_173_n374(net141_c1,net141);
INTERCONNECT Split_180_n381_NOTT_8_n44(net142_c1,net142);
INTERCONNECT Split_157_n358_OR2T_48_n84(net143_c1,net143);
INTERCONNECT Split_165_n366_OR2T_42_n78(net144_c1,net144);
INTERCONNECT Split_173_n374_AND2T_9_n45(net145_c1,net145);
INTERCONNECT Split_181_n382_Split_182_n383(net146_c1,net146);
INTERCONNECT Split_158_n359_OR2T_33_n69(net147_c1,net147);
INTERCONNECT Split_166_n367_DFFT_77__FBL_n278(net148_c1,net148);
INTERCONNECT Split_174_n375_AND2T_11_n47(net149_c1,net149);
INTERCONNECT Split_182_n383_NOTT_12_n48(net150_c1,net150);
INTERCONNECT Split_167_n368_OR2T_56_n92(net151_c1,net151);
INTERCONNECT Split_175_n376_DFFT_107__FPB_n308(net152_c1,net152);
INTERCONNECT Split_183_n384_XOR2T_29_n65(net153_c1,net153);
INTERCONNECT Split_168_n369_DFFT_78__FBL_n279(net154_c1,net154);
INTERCONNECT Split_176_n377_OR2T_49_n85(net155_c1,net155);
INTERCONNECT Split_184_n385_Split_185_n386(net156_c1,net156);
INTERCONNECT Split_177_n378_DFFT_120__FPB_n321(net157_c1,net157);
INTERCONNECT Split_185_n386_NOTT_13_n49(net158_c1,net158);
INTERCONNECT Split_178_n379_NOTT_15_n51(net159_c1,net159);
INTERCONNECT Split_186_n387_XOR2T_29_n65(net160_c1,net160);
INTERCONNECT DFFT_63_state_obs0_buf_DFFT_69__PIPL_n111(net161_c1,net161);
INTERCONNECT DFFT_64_state_obs1_buf_DFFT_70__PIPL_n112(net162_c1,net162);
INTERCONNECT DFFT_65_state_obs2_buf_DFFT_71__PIPL_n113(net163_c1,net163);
INTERCONNECT DFFT_66_state_obs3_buf_DFFT_72__PIPL_n114(net164_c1,net164);
INTERCONNECT DFFT_69__PIPL_n111_DFFT_121__FPB_n322(net165_c1,net165);
INTERCONNECT DFFT_70__PIPL_n112_DFFT_125__FPB_n326(net166_c1,net166);
INTERCONNECT DFFT_71__PIPL_n113_DFFT_129__FPB_n330(net167_c1,net167);
INTERCONNECT DFFT_72__PIPL_n114_DFFT_133__FPB_n334(net168_c1,net168);
INTERCONNECT DFFT_73__PIPL_n115_DFFT_63_state_obs0_buf(net169_c1,net169);
INTERCONNECT DFFT_74__PIPL_n116_DFFT_64_state_obs1_buf(net170_c1,net170);
INTERCONNECT DFFT_75__PIPL_n117_DFFT_65_state_obs2_buf(net171_c1,net171);
INTERCONNECT DFFT_76__PIPL_n118_DFFT_66_state_obs3_buf(net172_c1,net172);
INTERCONNECT DFFT_79__FBL_n280_Split_177_n378(net173_c1,net173);
INTERCONNECT DFFT_80__FBL_n281_Split_179_n380(net174_c1,net174);
INTERCONNECT DFFT_81__FBL_n282_Split_181_n382(net175_c1,net175);
INTERCONNECT DFFT_82__FBL_n283_Split_184_n385(net176_c1,net176);
INTERCONNECT DFFT_77__FBL_n278_DFFT_92__FPB_n293(net177_c1,net177);
INTERCONNECT DFFT_78__FBL_n279_Split_175_n376(net178_c1,net178);
INTERCONNECT DFFT_99__FPB_n300_DFFT_100__FPB_n301(net179_c1,net179);
INTERCONNECT DFFT_100__FPB_n301_DFFT_101__FPB_n302(net180_c1,net180);
INTERCONNECT DFFT_109__FPB_n310_DFFT_110__FPB_n311(net181_c1,net181);
INTERCONNECT DFFT_101__FPB_n302_OR2T_36_n72(net182_c1,net182);
INTERCONNECT DFFT_110__FPB_n311_DFFT_111__FPB_n312(net183_c1,net183);
INTERCONNECT DFFT_102__FPB_n303_AND2T_39_n75(net184_c1,net184);
INTERCONNECT DFFT_103__FPB_n304_DFFT_104__FPB_n305(net185_c1,net185);
INTERCONNECT DFFT_119__FPB_n320_AND2T_62_n98(net186_c1,net186);
INTERCONNECT DFFT_111__FPB_n312_AND2T_50_n86(net187_c1,net187);
INTERCONNECT DFFT_120__FPB_n321_AND2T_67_n109(net188_c1,net188);
INTERCONNECT DFFT_112__FPB_n313_OR2T_52_n88(net189_c1,net189);
INTERCONNECT DFFT_104__FPB_n305_OR2T_41_n77(net190_c1,net190);
INTERCONNECT DFFT_129__FPB_n330_DFFT_130__FPB_n331(net191_c1,net191);
INTERCONNECT DFFT_121__FPB_n322_DFFT_122__FPB_n323(net192_c1,net192);
INTERCONNECT DFFT_113__FPB_n314_DFFT_114__FPB_n315(net193_c1,net193);
INTERCONNECT DFFT_105__FPB_n306_AND2T_44_n80(net194_c1,net194);
INTERCONNECT DFFT_130__FPB_n331_DFFT_131__FPB_n332(net195_c1,net195);
INTERCONNECT DFFT_122__FPB_n323_DFFT_123__FPB_n324(net196_c1,net196);
INTERCONNECT DFFT_114__FPB_n315_AND2T_54_n90(net197_c1,net197);
INTERCONNECT DFFT_106__FPB_n307_AND2T_45_n81(net198_c1,net198);
INTERCONNECT DFFT_131__FPB_n332_DFFT_132_state_obs2(net199_c1,net199);
INTERCONNECT DFFT_123__FPB_n324_DFFT_124_state_obs0(net200_c1,net200);
INTERCONNECT DFFT_115__FPB_n316_AND2T_57_n93(net201_c1,net201);
INTERCONNECT DFFT_107__FPB_n308_AND2T_46_n82(net202_c1,net202);
INTERCONNECT DFFT_116__FPB_n317_AND2T_59_n95(net203_c1,net203);
INTERCONNECT DFFT_108__FPB_n309_AND2T_47_n83(net204_c1,net204);
INTERCONNECT DFFT_133__FPB_n334_DFFT_134__FPB_n335(net205_c1,net205);
INTERCONNECT DFFT_125__FPB_n326_DFFT_126__FPB_n327(net206_c1,net206);
INTERCONNECT DFFT_117__FPB_n318_AND2T_61_n97(net207_c1,net207);
INTERCONNECT DFFT_134__FPB_n335_DFFT_135_state_obs3(net208_c1,net208);
INTERCONNECT DFFT_126__FPB_n327_DFFT_127__FPB_n328(net209_c1,net209);
INTERCONNECT DFFT_118__FPB_n319_DFFT_119__FPB_n320(net210_c1,net210);
INTERCONNECT DFFT_127__FPB_n328_DFFT_128_state_obs1(net211_c1,net211);
INTERCONNECT DFFT_89__FPB_n290_AND2T_24_n60(net212_c1,net212);
INTERCONNECT DFFT_90__FPB_n291_AND2T_25_n61(net213_c1,net213);
INTERCONNECT DFFT_83__FPB_n284_DFFT_80__FBL_n281(net214_c1,net214);
INTERCONNECT DFFT_91__FPB_n292_AND2T_28_n64(net215_c1,net215);
INTERCONNECT DFFT_92__FPB_n293_AND2T_30_n66(net216_c1,net216);
INTERCONNECT DFFT_84__FPB_n285_AND2T_9_n45(net217_c1,net217);
INTERCONNECT DFFT_93__FPB_n294_OR2T_33_n69(net218_c1,net218);
INTERCONNECT DFFT_85__FPB_n286_AND2T_10_n46(net219_c1,net219);
INTERCONNECT DFFT_94__FPB_n295_DFFT_95__FPB_n296(net220_c1,net220);
INTERCONNECT DFFT_86__FPB_n287_AND2T_11_n47(net221_c1,net221);
INTERCONNECT DFFT_95__FPB_n296_DFFT_96__FPB_n297(net222_c1,net222);
INTERCONNECT DFFT_87__FPB_n288_AND2T_16_n52(net223_c1,net223);
INTERCONNECT DFFT_96__FPB_n297_DFFT_97__FPB_n298(net224_c1,net224);
INTERCONNECT DFFT_88__FPB_n289_AND2T_21_n57(net225_c1,net225);
INTERCONNECT DFFT_97__FPB_n298_DFFT_98__FPB_n299(net226_c1,net226);
INTERCONNECT DFFT_98__FPB_n299_AND2T_35_n71(net227_c1,net227);
INTERCONNECT DFFT_124_state_obs0_state_obs0_Pad(net228_c1,state_obs0_Pad);
INTERCONNECT DFFT_128_state_obs1_state_obs1_Pad(net229_c1,state_obs1_Pad);
INTERCONNECT DFFT_132_state_obs2_state_obs2_Pad(net230_c1,state_obs2_Pad);
INTERCONNECT DFFT_135_state_obs3_state_obs3_Pad(net231_c1,state_obs3_Pad);
INTERCONNECT SplitCLK_0_255_SplitCLK_0_191(net232_c1,net232);
INTERCONNECT SplitCLK_0_255_SplitCLK_2_254(net233_c1,net233);
INTERCONNECT SplitCLK_2_254_SplitCLK_6_222(net234_c1,net234);
INTERCONNECT SplitCLK_2_254_SplitCLK_4_253(net235_c1,net235);
INTERCONNECT SplitCLK_4_253_SplitCLK_4_237(net236_c1,net236);
INTERCONNECT SplitCLK_4_253_SplitCLK_2_252(net237_c1,net237);
INTERCONNECT SplitCLK_2_252_SplitCLK_6_244(net238_c1,net238);
INTERCONNECT SplitCLK_2_252_SplitCLK_4_251(net239_c1,net239);
INTERCONNECT SplitCLK_4_251_SplitCLK_0_247(net240_c1,net240);
INTERCONNECT SplitCLK_4_251_SplitCLK_6_250(net241_c1,net241);
INTERCONNECT SplitCLK_6_250_SplitCLK_0_248(net242_c1,net242);
INTERCONNECT SplitCLK_6_250_SplitCLK_4_249(net243_c1,net243);
INTERCONNECT SplitCLK_4_249_OR2T_49_n85(net244_c1,net244);
INTERCONNECT SplitCLK_4_249_DFFT_109__FPB_n310(net245_c1,net245);
INTERCONNECT SplitCLK_0_248_OR2T_52_n88(net246_c1,net246);
INTERCONNECT SplitCLK_0_248_DFFT_78__FBL_n279(net247_c1,net247);
INTERCONNECT SplitCLK_0_247_SplitCLK_0_245(net248_c1,net248);
INTERCONNECT SplitCLK_0_247_SplitCLK_4_246(net249_c1,net249);
INTERCONNECT SplitCLK_4_246_DFFT_99__FPB_n300(net250_c1,net250);
INTERCONNECT SplitCLK_4_246_DFFT_116__FPB_n317(net251_c1,net251);
INTERCONNECT SplitCLK_0_245_DFFT_110__FPB_n311(net252_c1,net252);
INTERCONNECT SplitCLK_0_245_DFFT_111__FPB_n312(net253_c1,net253);
INTERCONNECT SplitCLK_6_244_SplitCLK_0_240(net254_c1,net254);
INTERCONNECT SplitCLK_6_244_SplitCLK_2_243(net255_c1,net255);
INTERCONNECT SplitCLK_2_243_SplitCLK_4_241(net256_c1,net256);
INTERCONNECT SplitCLK_2_243_SplitCLK_4_242(net257_c1,net257);
INTERCONNECT SplitCLK_4_242_AND2T_43_n79(net258_c1,net258);
INTERCONNECT SplitCLK_4_242_AND2T_53_n89(net259_c1,net259);
INTERCONNECT SplitCLK_4_241_AND2T_44_n80(net260_c1,net260);
INTERCONNECT SplitCLK_4_241_DFFT_105__FPB_n306(net261_c1,net261);
INTERCONNECT SplitCLK_0_240_SplitCLK_4_238(net262_c1,net262);
INTERCONNECT SplitCLK_0_240_SplitCLK_4_239(net263_c1,net263);
INTERCONNECT SplitCLK_4_239_AND2T_51_n87(net264_c1,net264);
INTERCONNECT SplitCLK_4_239_DFFT_112__FPB_n313(net265_c1,net265);
INTERCONNECT SplitCLK_4_238_OR2T_33_n69(net266_c1,net266);
INTERCONNECT SplitCLK_4_238_DFFT_90__FPB_n291(net267_c1,net267);
INTERCONNECT SplitCLK_4_237_SplitCLK_6_229(net268_c1,net268);
INTERCONNECT SplitCLK_4_237_SplitCLK_4_236(net269_c1,net269);
INTERCONNECT SplitCLK_4_236_SplitCLK_4_232(net270_c1,net270);
INTERCONNECT SplitCLK_4_236_SplitCLK_2_235(net271_c1,net271);
INTERCONNECT SplitCLK_2_235_SplitCLK_4_233(net272_c1,net272);
INTERCONNECT SplitCLK_2_235_SplitCLK_4_234(net273_c1,net273);
INTERCONNECT SplitCLK_4_234_DFFT_100__FPB_n301(net274_c1,net274);
INTERCONNECT SplitCLK_4_234_DFFT_101__FPB_n302(net275_c1,net275);
INTERCONNECT SplitCLK_4_233_AND2T_50_n86(net276_c1,net276);
INTERCONNECT SplitCLK_4_233_OR2T_37_n73(net277_c1,net277);
INTERCONNECT SplitCLK_4_232_SplitCLK_4_230(net278_c1,net278);
INTERCONNECT SplitCLK_4_232_SplitCLK_4_231(net279_c1,net279);
INTERCONNECT SplitCLK_4_231_AND2T_59_n95(net280_c1,net280);
INTERCONNECT SplitCLK_4_231_NOTT_38_n74(net281_c1,net281);
INTERCONNECT SplitCLK_4_230_AND2T_39_n75(net282_c1,net282);
INTERCONNECT SplitCLK_4_230_DFFT_102__FPB_n303(net283_c1,net283);
INTERCONNECT SplitCLK_6_229_SplitCLK_0_225(net284_c1,net284);
INTERCONNECT SplitCLK_6_229_SplitCLK_6_228(net285_c1,net285);
INTERCONNECT SplitCLK_6_228_SplitCLK_4_226(net286_c1,net286);
INTERCONNECT SplitCLK_6_228_SplitCLK_4_227(net287_c1,net287);
INTERCONNECT SplitCLK_4_227_AND2T_45_n81(net288_c1,net288);
INTERCONNECT SplitCLK_4_227_DFFT_93__FPB_n294(net289_c1,net289);
INTERCONNECT SplitCLK_4_226_NOTT_58_n94(net290_c1,net290);
INTERCONNECT SplitCLK_4_226_DFFT_106__FPB_n307(net291_c1,net291);
INTERCONNECT SplitCLK_0_225_SplitCLK_0_223(net292_c1,net292);
INTERCONNECT SplitCLK_0_225_SplitCLK_4_224(net293_c1,net293);
INTERCONNECT SplitCLK_4_224_OR2T_42_n78(net294_c1,net294);
INTERCONNECT SplitCLK_4_224_OR2T_48_n84(net295_c1,net295);
INTERCONNECT SplitCLK_0_223_AND2T_25_n61(net296_c1,net296);
INTERCONNECT SplitCLK_0_223_DFFT_117__FPB_n318(net297_c1,net297);
INTERCONNECT SplitCLK_6_222_SplitCLK_6_206(net298_c1,net298);
INTERCONNECT SplitCLK_6_222_SplitCLK_6_221(net299_c1,net299);
INTERCONNECT SplitCLK_6_221_SplitCLK_6_213(net300_c1,net300);
INTERCONNECT SplitCLK_6_221_SplitCLK_6_220(net301_c1,net301);
INTERCONNECT SplitCLK_6_220_SplitCLK_0_216(net302_c1,net302);
INTERCONNECT SplitCLK_6_220_SplitCLK_2_219(net303_c1,net303);
INTERCONNECT SplitCLK_2_219_SplitCLK_4_217(net304_c1,net304);
INTERCONNECT SplitCLK_2_219_SplitCLK_4_218(net305_c1,net305);
INTERCONNECT SplitCLK_4_218_DFFT_81__FBL_n282(net306_c1,net306);
INTERCONNECT SplitCLK_4_218_DFFT_82__FBL_n283(net307_c1,net307);
INTERCONNECT SplitCLK_4_217_AND2T_20_n56(net308_c1,net308);
INTERCONNECT SplitCLK_4_217_DFFT_84__FPB_n285(net309_c1,net309);
INTERCONNECT SplitCLK_0_216_SplitCLK_4_214(net310_c1,net310);
INTERCONNECT SplitCLK_0_216_SplitCLK_4_215(net311_c1,net311);
INTERCONNECT SplitCLK_4_215_AND2T_19_n55(net312_c1,net312);
INTERCONNECT SplitCLK_4_215_NOTT_12_n48(net313_c1,net313);
INTERCONNECT SplitCLK_4_214_AND2T_9_n45(net314_c1,net314);
INTERCONNECT SplitCLK_4_214_AND2T_16_n52(net315_c1,net315);
INTERCONNECT SplitCLK_6_213_SplitCLK_4_209(net316_c1,net316);
INTERCONNECT SplitCLK_6_213_SplitCLK_6_212(net317_c1,net317);
INTERCONNECT SplitCLK_6_212_SplitCLK_0_210(net318_c1,net318);
INTERCONNECT SplitCLK_6_212_SplitCLK_4_211(net319_c1,net319);
INTERCONNECT SplitCLK_4_211_DFFT_121__FPB_n322(net320_c1,net320);
INTERCONNECT SplitCLK_4_211_DFFT_69__PIPL_n111(net321_c1,net321);
INTERCONNECT SplitCLK_0_210_DFFT_123__FPB_n324(net322_c1,net322);
INTERCONNECT SplitCLK_0_210_DFFT_124_state_obs0(net323_c1,net323);
INTERCONNECT SplitCLK_4_209_SplitCLK_0_207(net324_c1,net324);
INTERCONNECT SplitCLK_4_209_SplitCLK_4_208(net325_c1,net325);
INTERCONNECT SplitCLK_4_208_DFFT_63_state_obs0_buf(net326_c1,net326);
INTERCONNECT SplitCLK_4_208_DFFT_73__PIPL_n115(net327_c1,net327);
INTERCONNECT SplitCLK_0_207_DFFT_122__FPB_n323(net328_c1,net328);
INTERCONNECT SplitCLK_0_207_DFFT_128_state_obs1(net329_c1,net329);
INTERCONNECT SplitCLK_6_206_SplitCLK_6_198(net330_c1,net330);
INTERCONNECT SplitCLK_6_206_SplitCLK_4_205(net331_c1,net331);
INTERCONNECT SplitCLK_4_205_SplitCLK_4_201(net332_c1,net332);
INTERCONNECT SplitCLK_4_205_SplitCLK_6_204(net333_c1,net333);
INTERCONNECT SplitCLK_6_204_SplitCLK_0_202(net334_c1,net334);
INTERCONNECT SplitCLK_6_204_SplitCLK_4_203(net335_c1,net335);
INTERCONNECT SplitCLK_4_203_AND2T_11_n47(net336_c1,net336);
INTERCONNECT SplitCLK_4_203_DFFT_77__FBL_n278(net337_c1,net337);
INTERCONNECT SplitCLK_0_202_AND2T_10_n46(net338_c1,net338);
INTERCONNECT SplitCLK_0_202_DFFT_85__FPB_n286(net339_c1,net339);
INTERCONNECT SplitCLK_4_201_SplitCLK_4_199(net340_c1,net340);
INTERCONNECT SplitCLK_4_201_SplitCLK_4_200(net341_c1,net341);
INTERCONNECT SplitCLK_4_200_NOTT_13_n49(net342_c1,net342);
INTERCONNECT SplitCLK_4_200_DFFT_92__FPB_n293(net343_c1,net343);
INTERCONNECT SplitCLK_4_199_XOR2T_29_n65(net344_c1,net344);
INTERCONNECT SplitCLK_4_199_AND2T_17_n53(net345_c1,net345);
INTERCONNECT SplitCLK_6_198_SplitCLK_4_194(net346_c1,net346);
INTERCONNECT SplitCLK_6_198_SplitCLK_6_197(net347_c1,net347);
INTERCONNECT SplitCLK_6_197_SplitCLK_0_195(net348_c1,net348);
INTERCONNECT SplitCLK_6_197_SplitCLK_4_196(net349_c1,net349);
INTERCONNECT SplitCLK_4_196_DFFT_64_state_obs1_buf(net350_c1,net350);
INTERCONNECT SplitCLK_4_196_DFFT_74__PIPL_n116(net351_c1,net351);
INTERCONNECT SplitCLK_0_195_DFFT_126__FPB_n327(net352_c1,net352);
INTERCONNECT SplitCLK_0_195_DFFT_127__FPB_n328(net353_c1,net353);
INTERCONNECT SplitCLK_4_194_SplitCLK_0_192(net354_c1,net354);
INTERCONNECT SplitCLK_4_194_SplitCLK_4_193(net355_c1,net355);
INTERCONNECT SplitCLK_4_193_DFFT_70__PIPL_n112(net356_c1,net356);
INTERCONNECT SplitCLK_4_193_DFFT_125__FPB_n326(net357_c1,net357);
INTERCONNECT SplitCLK_0_192_DFFT_131__FPB_n332(net358_c1,net358);
INTERCONNECT SplitCLK_0_192_DFFT_132_state_obs2(net359_c1,net359);
INTERCONNECT SplitCLK_0_191_SplitCLK_6_159(net360_c1,net360);
INTERCONNECT SplitCLK_0_191_SplitCLK_4_190(net361_c1,net361);
INTERCONNECT SplitCLK_4_190_SplitCLK_0_174(net362_c1,net362);
INTERCONNECT SplitCLK_4_190_SplitCLK_4_189(net363_c1,net363);
INTERCONNECT SplitCLK_4_189_SplitCLK_2_181(net364_c1,net364);
INTERCONNECT SplitCLK_4_189_SplitCLK_4_188(net365_c1,net365);
INTERCONNECT SplitCLK_4_188_SplitCLK_0_184(net366_c1,net366);
INTERCONNECT SplitCLK_4_188_SplitCLK_6_187(net367_c1,net367);
INTERCONNECT SplitCLK_6_187_SplitCLK_4_185(net368_c1,net368);
INTERCONNECT SplitCLK_6_187_SplitCLK_4_186(net369_c1,net369);
INTERCONNECT SplitCLK_4_186_OR2T_36_n72(net370_c1,net370);
INTERCONNECT SplitCLK_4_186_DFFT_96__FPB_n297(net371_c1,net371);
INTERCONNECT SplitCLK_4_185_AND2T_40_n76(net372_c1,net372);
INTERCONNECT SplitCLK_4_185_DFFT_107__FPB_n308(net373_c1,net373);
INTERCONNECT SplitCLK_0_184_SplitCLK_4_182(net374_c1,net374);
INTERCONNECT SplitCLK_0_184_SplitCLK_4_183(net375_c1,net375);
INTERCONNECT SplitCLK_4_183_DFFT_97__FPB_n298(net376_c1,net376);
INTERCONNECT SplitCLK_4_183_DFFT_98__FPB_n299(net377_c1,net377);
INTERCONNECT SplitCLK_4_182_AND2T_46_n82(net378_c1,net378);
INTERCONNECT SplitCLK_4_182_DFFT_108__FPB_n309(net379_c1,net379);
INTERCONNECT SplitCLK_2_181_SplitCLK_4_177(net380_c1,net380);
INTERCONNECT SplitCLK_2_181_SplitCLK_6_180(net381_c1,net381);
INTERCONNECT SplitCLK_6_180_SplitCLK_0_178(net382_c1,net382);
INTERCONNECT SplitCLK_6_180_SplitCLK_4_179(net383_c1,net383);
INTERCONNECT SplitCLK_4_179_AND2T_60_n96(net384_c1,net384);
INTERCONNECT SplitCLK_4_179_AND2T_61_n97(net385_c1,net385);
INTERCONNECT SplitCLK_0_178_DFFT_118__FPB_n319(net386_c1,net386);
INTERCONNECT SplitCLK_0_178_DFFT_119__FPB_n320(net387_c1,net387);
INTERCONNECT SplitCLK_4_177_SplitCLK_0_175(net388_c1,net388);
INTERCONNECT SplitCLK_4_177_SplitCLK_4_176(net389_c1,net389);
INTERCONNECT SplitCLK_4_176_AND2T_47_n83(net390_c1,net390);
INTERCONNECT SplitCLK_4_176_OR2T_41_n77(net391_c1,net391);
INTERCONNECT SplitCLK_0_175_OR2T_34_n70(net392_c1,net392);
INTERCONNECT SplitCLK_0_175_OR2T_27_n63(net393_c1,net393);
INTERCONNECT SplitCLK_0_174_SplitCLK_4_166(net394_c1,net394);
INTERCONNECT SplitCLK_0_174_SplitCLK_4_173(net395_c1,net395);
INTERCONNECT SplitCLK_4_173_SplitCLK_0_169(net396_c1,net396);
INTERCONNECT SplitCLK_4_173_SplitCLK_4_172(net397_c1,net397);
INTERCONNECT SplitCLK_4_172_SplitCLK_4_170(net398_c1,net398);
INTERCONNECT SplitCLK_4_172_SplitCLK_4_171(net399_c1,net399);
INTERCONNECT SplitCLK_4_171_DFFT_94__FPB_n295(net400_c1,net400);
INTERCONNECT SplitCLK_4_171_DFFT_95__FPB_n296(net401_c1,net401);
INTERCONNECT SplitCLK_4_170_NOTT_18_n54(net402_c1,net402);
INTERCONNECT SplitCLK_4_170_DFFT_103__FPB_n304(net403_c1,net403);
INTERCONNECT SplitCLK_0_169_SplitCLK_0_167(net404_c1,net404);
INTERCONNECT SplitCLK_0_169_SplitCLK_4_168(net405_c1,net405);
INTERCONNECT SplitCLK_4_168_DFFT_113__FPB_n314(net406_c1,net406);
INTERCONNECT SplitCLK_4_168_DFFT_114__FPB_n315(net407_c1,net407);
INTERCONNECT SplitCLK_0_167_OR2T_26_n62(net408_c1,net408);
INTERCONNECT SplitCLK_0_167_DFFT_104__FPB_n305(net409_c1,net409);
INTERCONNECT SplitCLK_4_166_SplitCLK_0_162(net410_c1,net410);
INTERCONNECT SplitCLK_4_166_SplitCLK_6_165(net411_c1,net411);
INTERCONNECT SplitCLK_6_165_SplitCLK_0_163(net412_c1,net412);
INTERCONNECT SplitCLK_6_165_SplitCLK_4_164(net413_c1,net413);
INTERCONNECT SplitCLK_4_164_AND2T_35_n71(net414_c1,net414);
INTERCONNECT SplitCLK_4_164_OR2T_55_n91(net415_c1,net415);
INTERCONNECT SplitCLK_0_163_AND2T_62_n98(net416_c1,net416);
INTERCONNECT SplitCLK_0_163_AND2T_57_n93(net417_c1,net417);
INTERCONNECT SplitCLK_0_162_SplitCLK_0_160(net418_c1,net418);
INTERCONNECT SplitCLK_0_162_SplitCLK_4_161(net419_c1,net419);
INTERCONNECT SplitCLK_4_161_AND2T_54_n90(net420_c1,net420);
INTERCONNECT SplitCLK_4_161_OR2T_56_n92(net421_c1,net421);
INTERCONNECT SplitCLK_0_160_DFFT_115__FPB_n316(net422_c1,net422);
INTERCONNECT SplitCLK_0_160_DFFT_79__FBL_n280(net423_c1,net423);
INTERCONNECT SplitCLK_6_159_SplitCLK_0_143(net424_c1,net424);
INTERCONNECT SplitCLK_6_159_SplitCLK_2_158(net425_c1,net425);
INTERCONNECT SplitCLK_2_158_SplitCLK_6_150(net426_c1,net426);
INTERCONNECT SplitCLK_2_158_SplitCLK_4_157(net427_c1,net427);
INTERCONNECT SplitCLK_4_157_SplitCLK_4_153(net428_c1,net428);
INTERCONNECT SplitCLK_4_157_SplitCLK_6_156(net429_c1,net429);
INTERCONNECT SplitCLK_6_156_SplitCLK_4_154(net430_c1,net430);
INTERCONNECT SplitCLK_6_156_SplitCLK_4_155(net431_c1,net431);
INTERCONNECT SplitCLK_4_155_AND2T_21_n57(net432_c1,net432);
INTERCONNECT SplitCLK_4_155_OR2T_32_n68(net433_c1,net433);
INTERCONNECT SplitCLK_4_154_AND2T_31_n67(net434_c1,net434);
INTERCONNECT SplitCLK_4_154_NOTT_15_n51(net435_c1,net435);
INTERCONNECT SplitCLK_4_153_SplitCLK_4_151(net436_c1,net436);
INTERCONNECT SplitCLK_4_153_SplitCLK_4_152(net437_c1,net437);
INTERCONNECT SplitCLK_4_152_OR2T_23_n59(net438_c1,net438);
INTERCONNECT SplitCLK_4_152_DFFT_88__FPB_n289(net439_c1,net439);
INTERCONNECT SplitCLK_4_151_AND2T_30_n66(net440_c1,net440);
INTERCONNECT SplitCLK_4_151_DFFT_86__FPB_n287(net441_c1,net441);
INTERCONNECT SplitCLK_6_150_SplitCLK_2_146(net442_c1,net442);
INTERCONNECT SplitCLK_6_150_SplitCLK_2_149(net443_c1,net443);
INTERCONNECT SplitCLK_2_149_SplitCLK_4_147(net444_c1,net444);
INTERCONNECT SplitCLK_2_149_SplitCLK_4_148(net445_c1,net445);
INTERCONNECT SplitCLK_4_148_AND2T_28_n64(net446_c1,net446);
INTERCONNECT SplitCLK_4_148_DFFT_91__FPB_n292(net447_c1,net447);
INTERCONNECT SplitCLK_4_147_DFFT_65_state_obs2_buf(net448_c1,net448);
INTERCONNECT SplitCLK_4_147_DFFT_130__FPB_n331(net449_c1,net449);
INTERCONNECT SplitCLK_2_146_SplitCLK_4_144(net450_c1,net450);
INTERCONNECT SplitCLK_2_146_SplitCLK_4_145(net451_c1,net451);
INTERCONNECT SplitCLK_4_145_DFFT_71__PIPL_n113(net452_c1,net452);
INTERCONNECT SplitCLK_4_145_DFFT_75__PIPL_n117(net453_c1,net453);
INTERCONNECT SplitCLK_4_144_DFFT_129__FPB_n330(net454_c1,net454);
INTERCONNECT SplitCLK_4_144_DFFT_135_state_obs3(net455_c1,net455);
INTERCONNECT SplitCLK_0_143_SplitCLK_6_135(net456_c1,net456);
INTERCONNECT SplitCLK_0_143_SplitCLK_4_142(net457_c1,net457);
INTERCONNECT SplitCLK_4_142_SplitCLK_0_138(net458_c1,net458);
INTERCONNECT SplitCLK_4_142_SplitCLK_2_141(net459_c1,net459);
INTERCONNECT SplitCLK_2_141_SplitCLK_0_139(net460_c1,net460);
INTERCONNECT SplitCLK_2_141_SplitCLK_4_140(net461_c1,net461);
INTERCONNECT SplitCLK_4_140_AND2T_14_n50(net462_c1,net462);
INTERCONNECT SplitCLK_4_140_DFFT_89__FPB_n290(net463_c1,net463);
INTERCONNECT SplitCLK_0_139_DFFT_120__FPB_n321(net464_c1,net464);
INTERCONNECT SplitCLK_0_139_DFFT_87__FPB_n288(net465_c1,net465);
INTERCONNECT SplitCLK_0_138_SplitCLK_4_136(net466_c1,net466);
INTERCONNECT SplitCLK_0_138_SplitCLK_4_137(net467_c1,net467);
INTERCONNECT SplitCLK_4_137_AND2T_24_n60(net468_c1,net468);
INTERCONNECT SplitCLK_4_137_DFFT_83__FPB_n284(net469_c1,net469);
INTERCONNECT SplitCLK_4_136_AND2T_22_n58(net470_c1,net470);
INTERCONNECT SplitCLK_4_136_DFFT_80__FBL_n281(net471_c1,net471);
INTERCONNECT SplitCLK_6_135_SplitCLK_4_131(net472_c1,net472);
INTERCONNECT SplitCLK_6_135_SplitCLK_2_134(net473_c1,net473);
INTERCONNECT SplitCLK_2_134_SplitCLK_4_132(net474_c1,net474);
INTERCONNECT SplitCLK_2_134_SplitCLK_4_133(net475_c1,net475);
INTERCONNECT SplitCLK_4_133_NOTT_8_n44(net476_c1,net476);
INTERCONNECT SplitCLK_4_133_AND2T_67_n109(net477_c1,net477);
INTERCONNECT SplitCLK_4_132_DFFT_66_state_obs3_buf(net478_c1,net478);
INTERCONNECT SplitCLK_4_132_DFFT_76__PIPL_n118(net479_c1,net479);
INTERCONNECT SplitCLK_4_131_SplitCLK_4_129(net480_c1,net480);
INTERCONNECT SplitCLK_4_131_SplitCLK_4_130(net481_c1,net481);
INTERCONNECT SplitCLK_4_130_DFFT_72__PIPL_n114(net482_c1,net482);
INTERCONNECT SplitCLK_4_130_NOTT_68_n110(net483_c1,net483);
INTERCONNECT SplitCLK_4_129_DFFT_133__FPB_n334(net484_c1,net484);
INTERCONNECT SplitCLK_4_129_DFFT_134__FPB_n335(net485_c1,net485);
INTERCONNECT GCLK_Pad_SplitCLK_0_255(GCLK_Pad,net486);

endmodule
