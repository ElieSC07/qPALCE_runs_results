module TAP_half_route(
input GCLK_Pad,
input TMS_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output state_obs2_Pad,
output state_obs3_Pad);

wire TMS_Pad;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire TRST_Pad;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire state_obs0_Pad;
wire net229_c1;
wire state_obs1_Pad;
wire net230_c1;
wire state_obs2_Pad;
wire net231_c1;
wire state_obs3_Pad;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire GCLK_Pad;
wire net486;

DFFT DFFT_99__FPB_n312(net372,net155,net175_c1);
XOR2T XOR2T_29_n53(net344,net160,net156,net16_c1);
AND2T AND2T_9_n33(net314,net150,net221,net4_c1);
NOTT NOTT_8_n32(net476,net148,net2_c1);
AND2T AND2T_10_n34(net315,net99,net210,net7_c1);
AND2T AND2T_11_n35(net432,net153,net213,net10_c1);
AND2T AND2T_20_n44(net338,net103,net83,net13_c1);
AND2T AND2T_21_n45(net296,net121,net215,net17_c1);
AND2T AND2T_30_n54(net440,net73,net220,net21_c1);
AND2T AND2T_22_n46(net470,net78,net140,net22_c1);
AND2T AND2T_14_n38(net312,net124,net118,net23_c1);
AND2T AND2T_31_n55(net441,net21,net116,net26_c1);
AND2T AND2T_16_n40(net313,net133,net214,net1_c1);
AND2T AND2T_40_n64(net408,net25,net112,net31_c1);
AND2T AND2T_24_n48(net438,net87,net216,net33_c1);
AND2T AND2T_17_n41(net345,net1,net128,net3_c1);
AND2T AND2T_25_n49(net439,net69,net217,net38_c1);
AND2T AND2T_50_n74(net276,net85,net190,net40_c1);
AND2T AND2T_19_n43(net306,net108,net102,net9_c1);
AND2T AND2T_51_n75(net264,net40,net30,net44_c1);
AND2T AND2T_43_n67(net265,net41,net15,net45_c1);
AND2T AND2T_35_n59(net390,net122,net172,net46_c1);
AND2T AND2T_28_n52(net446,net144,net219,net12_c1);
AND2T AND2T_60_n84(net422,net43,net61,net47_c1);
AND2T AND2T_44_n68(net258,net135,net170,net49_c1);
AND2T AND2T_61_n85(net414,net47,net181,net51_c1);
AND2T AND2T_53_n77(net259,net48,net81,net52_c1);
AND2T AND2T_45_n69(net288,net98,net171,net53_c1);
AND2T AND2T_46_n70(net378,net146,net175,net19_c1);
AND2T AND2T_62_n86(net423,net72,net189,net55_c1);
AND2T AND2T_54_n78(net409,net82,net202,net56_c1);
AND2T AND2T_47_n71(net384,net138,net178,net24_c1);
AND2T AND2T_39_n63(net289,net66,net185,net25_c1);
AND2T AND2T_63_n93(net477,net2,net193,net50_c1);
AND2T AND2T_57_n81(net386,net130,net174,net34_c1);
AND2T AND2T_59_n83(net406,net113,net177,net43_c1);
OR2T OR2T_23_n47(net387,net22,net17,net27_c1);
OR2T OR2T_32_n56(net433,net26,net137,net32_c1);
OR2T OR2T_41_n65(net420,net31,net195,net36_c1);
OR2T OR2T_33_n57(net266,net119,net222,net37_c1);
OR2T OR2T_26_n50(net402,net142,net134,net5_c1);
OR2T OR2T_42_n66(net294,net149,net77,net41_c1);
OR2T OR2T_34_n58(net392,net37,net8,net42_c1);
OR2T OR2T_27_n51(net415,net5,net129,net8_c1);
OR2T OR2T_36_n60(net373,net92,net182,net11_c1);
OR2T OR2T_52_n76(net246,net44,net194,net48_c1);
OR2T OR2T_37_n61(net277,net139,net68,net15_c1);
OR2T OR2T_55_n79(net391,net56,net125,net57_c1);
OR2T OR2T_56_n80(net385,net57,net123,net29_c1);
OR2T OR2T_48_n72(net295,net24,net117,net30_c1);
OR2T OR2T_49_n73(net244,net157,net58,net35_c1);
NOTT NOTT_12_n36(net260,net154,net14_c1);
NOTT NOTT_13_n37(net336,net159,net18_c1);
NOTT NOTT_15_n39(net308,net136,net28_c1);
NOTT NOTT_18_n42(net400,net100,net6_c1);
NOTT NOTT_38_n62(net280,net110,net20_c1);
NOTT NOTT_64_n94(net482,net96,net54_c1);
NOTT NOTT_58_n82(net468,net120,net39_c1);
DFFT DFFT_100__FPB_n313(net379,net19,net178_c1);
DFFT DFFT_101__FPB_n314(net245,net35,net180_c1);
DFFT DFFT_110__FPB_n323(net416,net51,net183_c1);
DFFT DFFT_102__FPB_n315(net250,net180,net184_c1);
DFFT DFFT_111__FPB_n324(net417,net183,net189_c1);
DFFT DFFT_103__FPB_n316(net252,net184,net190_c1);
DFFT DFFT_120__FPB_n333(net356,net187,net192_c1);
DFFT DFFT_112__FPB_n325(net464,net132,net193_c1);
DFFT DFFT_104__FPB_n317(net253,net70,net194_c1);
DFFT DFFT_121__FPB_n334(net357,net192,net197_c1);
DFFT DFFT_113__FPB_n326(net326,net224,net198_c1);
DFFT DFFT_105__FPB_n318(net403,net143,net199_c1);
DFFT DFFT_122__FPB_n335(net352,net197,net200_c1);
DFFT DFFT_114__FPB_n327(net320,net198,net201_c1);
DFFT DFFT_106__FPB_n319(net401,net199,net202_c1);
DFFT DFFT_107__FPB_n320(net297,net29,net174_c1);
DFFT DFFT_131__FPB_n344(net478,net227,net203_c1);
DFFT DFFT_123__FPB_n336(net353,net200,net204_c1);
DFFT DFFT_115__FPB_n328(net321,net201,net205_c1);
DFFT DFFT_108__FPB_n321(net251,net59,net177_c1);
DFFT DFFT_132__FPB_n345(net479,net203,net206_c1);
DFFT DFFT_116__FPB_n329(net328,net205,net207_c1);
DFFT DFFT_117__FPB_n330(net322,net207,net179_c1);
DFFT DFFT_109__FPB_n322(net393,net39,net181_c1);
DFFT DFFT_133__FPB_n346(net484,net206,net208_c1);
DFFT DFFT_125__FPB_n338(net447,net226,net209_c1);
DFFT DFFT_134__FPB_n347(net485,net208,net211_c1);
DFFT DFFT_126__FPB_n339(net452,net209,net212_c1);
DFFT DFFT_127__FPB_n340(net453,net212,net186_c1);
DFFT DFFT_119__FPB_n332(net350,net225,net187_c1);
DFFT DFFT_128__FPB_n341(net448,net186,net191_c1);
DFFT DFFT_129__FPB_n342(net358,net191,net196_c1);
DFFT DFFT_130_state_obs2(net359,net196,net230_c1);
DFFT DFFT_70__FBL_n283(net247,net126,net162_c1);
DFFT DFFT_71__FBL_n284(net462,net34,net163_c1);
DFFT DFFT_72__FBL_n285(net483,net218,net164_c1);
DFFT DFFT_80__FPB_n293(net342,net114,net215_c1);
DFFT DFFT_73__FBL_n286(net307,net101,net165_c1);
DFFT DFFT_81__FPB_n294(net337,net63,net216_c1);
DFFT DFFT_124_state_obs1(net329,net204,net229_c1);
DFFT DFFT_74__FBL_n287(net267,net75,net166_c1);
DFFT DFFT_90__FPB_n303(net370,net169,net172_c1);
DFFT DFFT_82__FPB_n295(net463,net67,net217_c1);
DFFT DFFT_65__PIPL_n95(net327,net4,net224_c1);
SPLITT Split_140_n353(net14,net62_c1,net115_c1);
SPLITT Split_141_n354(net115,net66_c1,net118_c1);
SPLITT Split_142_n355(net62,net67_c1,net120_c1);
SPLITT Split_150_n363(net65,net69_c1,net121_c1);
SPLITT Split_143_n356(net18,net73_c1,net124_c1);
SPLITT Split_151_n364(net27,net71_c1,net125_c1);
SPLITT Split_136_n349(net0,net74_c1,net127_c1);
SPLITT Split_144_n357(net23,net78_c1,net128_c1);
SPLITT Split_152_n365(net71,net77_c1,net129_c1);
SPLITT Split_160_n373(net46,net76_c1,net130_c1);
SPLITT Split_137_n350(net127,net58_c1,net110_c1);
SPLITT Split_145_n358(net28,net83_c1,net133_c1);
SPLITT Split_153_n366(net33,net82_c1,net134_c1);
SPLITT Split_161_n374(net76,net81_c1,net135_c1);
SPLITT Split_138_n351(net74,net59_c1,net111_c1);
SPLITT Split_146_n359(net3,net86_c1,net137_c1);
SPLITT Split_154_n367(net38,net84_c1,net138_c1);
SPLITT Split_162_n375(net11,net85_c1,net139_c1);
SPLITT Split_170_n383(net131,net87_c1,net140_c1);
SPLITT Split_139_n352(net10,net61_c1,net112_c1);
SPLITT Split_147_n360(net6,net60_c1,net113_c1);
SPLITT Split_155_n368(net84,net92_c1,net142_c1);
SPLITT Split_163_n376(net20,net89_c1,net143_c1);
SPLITT Split_171_n384(net79,net91_c1,net144_c1);
SPLITT Split_148_n361(net9,net63_c1,net114_c1);
SPLITT Split_156_n369(net12,net94_c1,net145_c1);
SPLITT Split_164_n377(net89,net95_c1,net146_c1);
SPLITT Split_172_n385(net54,net93_c1,net147_c1);
SPLITT Split_180_n393(net90,net96_c1,net148_c1);
SPLITT Split_149_n362(net13,net65_c1,net116_c1);
SPLITT Split_157_n370(net32,net64_c1,net117_c1);
SPLITT Split_165_n378(net36,net98_c1,net149_c1);
SPLITT Split_173_n386(net147,net99_c1,net150_c1);
SPLITT Split_181_n394(net165,net97_c1,net151_c1);
SPLITT Split_158_n371(net64,net68_c1,net119_c1);
SPLITT Split_166_n379(net49,net101_c1,net152_c1);
SPLITT Split_174_n387(net93,net103_c1,net153_c1);
SPLITT Split_182_n395(net151,net102_c1,net154_c1);
SPLITT Split_159_n372(net42,net72_c1,net122_c1);
SPLITT Split_167_n380(net53,net70_c1,net123_c1);
SPLITT Split_175_n388(net162,net104_c1,net155_c1);
SPLITT Split_183_n396(net97,net105_c1,net156_c1);
SPLITT Split_168_n381(net52,net75_c1,net126_c1);
SPLITT Split_176_n389(net104,net107_c1,net157_c1);
SPLITT Split_184_n397(net166,net106_c1,net158_c1);
SPLITT Split_169_n382(net50,net79_c1,net131_c1);
SPLITT Split_177_n390(net163,net80_c1,net132_c1);
SPLITT Split_185_n398(net158,net108_c1,net159_c1);
DFFT DFFT_91__FPB_n304(net274,net111,net173_c1);
SPLITT Split_178_n391(net80,net88_c1,net136_c1);
DFFT DFFT_83__FPB_n296(net434,net16,net219_c1);
DFFT DFFT_75__FPB_n288(net469,net55,net218_c1);
SPLITT Split_186_n399(net106,net109_c1,net160_c1);
SPLITT Split_179_n392(net164,net90_c1,net141_c1);
DFFT DFFT_66__PIPL_n96(net351,net7,net225_c1);
DFFT DFFT_92__FPB_n305(net275,net173,net176_c1);
DFFT DFFT_84__FPB_n297(net465,net161,net220_c1);
DFFT DFFT_76__FPB_n289(net309,net105,net221_c1);
DFFT DFFT_67__PIPL_n97(net449,net91,net226_c1);
DFFT DFFT_69__FBL_n282(net343,net152,net161_c1);
DFFT DFFT_93__FPB_n306(net281,net176,net182_c1);
DFFT DFFT_77__FPB_n290(net339,net109,net210_c1);
DFFT DFFT_85__FPB_n298(net290,net145,net222_c1);
DFFT DFFT_68__PIPL_n98(net454,net86,net227_c1);
DFFT DFFT_118_state_obs0(net323,net179,net228_c1);
DFFT DFFT_94__FPB_n307(net282,net107,net185_c1);
DFFT DFFT_78__FPB_n291(net435,net88,net213_c1);
DFFT DFFT_86__FPB_n299(net376,net60,net223_c1);
DFFT DFFT_87__FPB_n300(net377,net223,net167_c1);
DFFT DFFT_95__FPB_n308(net407,net95,net188_c1);
DFFT DFFT_79__FPB_n292(net471,net141,net214_c1);
DFFT DFFT_135_state_obs3(net455,net211,net231_c1);
DFFT DFFT_88__FPB_n301(net371,net167,net168_c1);
DFFT DFFT_96__FPB_n309(net421,net188,net195_c1);
DFFT DFFT_97__FPB_n310(net261,net45,net170_c1);
DFFT DFFT_89__FPB_n302(net283,net168,net169_c1);
DFFT DFFT_98__FPB_n311(net291,net94,net171_c1);
SPLITT SplitCLK_0_129(net480,net484_c1,net485_c1);
SPLITT SplitCLK_4_130(net481,net482_c1,net483_c1);
SPLITT SplitCLK_4_131(net472,net481_c1,net480_c1);
SPLITT SplitCLK_0_132(net474,net478_c1,net479_c1);
SPLITT SplitCLK_4_133(net475,net477_c1,net476_c1);
SPLITT SplitCLK_6_134(net473,net474_c1,net475_c1);
SPLITT SplitCLK_6_135(net456,net472_c1,net473_c1);
SPLITT SplitCLK_4_136(net466,net471_c1,net470_c1);
SPLITT SplitCLK_4_137(net467,net468_c1,net469_c1);
SPLITT SplitCLK_4_138(net458,net466_c1,net467_c1);
SPLITT SplitCLK_4_139(net460,net465_c1,net464_c1);
SPLITT SplitCLK_4_140(net461,net462_c1,net463_c1);
SPLITT SplitCLK_2_141(net459,net461_c1,net460_c1);
SPLITT SplitCLK_4_142(net457,net459_c1,net458_c1);
SPLITT SplitCLK_0_143(net424,net456_c1,net457_c1);
SPLITT SplitCLK_4_144(net450,net455_c1,net454_c1);
SPLITT SplitCLK_4_145(net451,net452_c1,net453_c1);
SPLITT SplitCLK_4_146(net442,net450_c1,net451_c1);
SPLITT SplitCLK_4_147(net444,net448_c1,net449_c1);
SPLITT SplitCLK_4_148(net445,net447_c1,net446_c1);
SPLITT SplitCLK_6_149(net443,net445_c1,net444_c1);
SPLITT SplitCLK_6_150(net426,net442_c1,net443_c1);
SPLITT SplitCLK_0_151(net436,net440_c1,net441_c1);
SPLITT SplitCLK_4_152(net437,net438_c1,net439_c1);
SPLITT SplitCLK_4_153(net428,net436_c1,net437_c1);
SPLITT SplitCLK_4_154(net430,net434_c1,net435_c1);
SPLITT SplitCLK_4_155(net431,net433_c1,net432_c1);
SPLITT SplitCLK_2_156(net429,net430_c1,net431_c1);
SPLITT SplitCLK_4_157(net427,net429_c1,net428_c1);
SPLITT SplitCLK_6_158(net425,net427_c1,net426_c1);
SPLITT SplitCLK_6_159(net360,net424_c1,net425_c1);
SPLITT SplitCLK_4_160(net418,net422_c1,net423_c1);
SPLITT SplitCLK_4_161(net419,net420_c1,net421_c1);
SPLITT SplitCLK_4_162(net410,net418_c1,net419_c1);
SPLITT SplitCLK_4_163(net412,net416_c1,net417_c1);
SPLITT SplitCLK_4_164(net413,net414_c1,net415_c1);
SPLITT SplitCLK_6_165(net411,net412_c1,net413_c1);
SPLITT SplitCLK_0_166(net394,net411_c1,net410_c1);
SPLITT SplitCLK_0_167(net404,net408_c1,net409_c1);
SPLITT SplitCLK_4_168(net405,net406_c1,net407_c1);
SPLITT SplitCLK_0_169(net396,net404_c1,net405_c1);
SPLITT SplitCLK_4_170(net398,net402_c1,net403_c1);
SPLITT SplitCLK_4_171(net399,net400_c1,net401_c1);
SPLITT SplitCLK_2_172(net397,net398_c1,net399_c1);
SPLITT SplitCLK_4_173(net395,net397_c1,net396_c1);
SPLITT SplitCLK_0_174(net362,net394_c1,net395_c1);
SPLITT SplitCLK_4_175(net388,net393_c1,net392_c1);
SPLITT SplitCLK_4_176(net389,net391_c1,net390_c1);
SPLITT SplitCLK_4_177(net380,net389_c1,net388_c1);
SPLITT SplitCLK_4_178(net382,net387_c1,net386_c1);
SPLITT SplitCLK_4_179(net383,net385_c1,net384_c1);
SPLITT SplitCLK_2_180(net381,net383_c1,net382_c1);
SPLITT SplitCLK_2_181(net364,net380_c1,net381_c1);
SPLITT SplitCLK_0_182(net374,net378_c1,net379_c1);
SPLITT SplitCLK_4_183(net375,net377_c1,net376_c1);
SPLITT SplitCLK_0_184(net366,net374_c1,net375_c1);
SPLITT SplitCLK_4_185(net368,net373_c1,net372_c1);
SPLITT SplitCLK_4_186(net369,net370_c1,net371_c1);
SPLITT SplitCLK_2_187(net367,net369_c1,net368_c1);
SPLITT SplitCLK_4_188(net365,net367_c1,net366_c1);
SPLITT SplitCLK_2_189(net363,net365_c1,net364_c1);
SPLITT SplitCLK_4_190(net361,net363_c1,net362_c1);
SPLITT SplitCLK_0_191(net232,net360_c1,net361_c1);
SPLITT SplitCLK_0_192(net354,net358_c1,net359_c1);
SPLITT SplitCLK_4_193(net355,net356_c1,net357_c1);
SPLITT SplitCLK_4_194(net346,net354_c1,net355_c1);
SPLITT SplitCLK_0_195(net348,net352_c1,net353_c1);
SPLITT SplitCLK_4_196(net349,net351_c1,net350_c1);
SPLITT SplitCLK_6_197(net347,net348_c1,net349_c1);
SPLITT SplitCLK_6_198(net330,net346_c1,net347_c1);
SPLITT SplitCLK_4_199(net340,net344_c1,net345_c1);
SPLITT SplitCLK_4_200(net341,net343_c1,net342_c1);
SPLITT SplitCLK_0_201(net332,net340_c1,net341_c1);
SPLITT SplitCLK_4_202(net334,net338_c1,net339_c1);
SPLITT SplitCLK_4_203(net335,net336_c1,net337_c1);
SPLITT SplitCLK_2_204(net333,net335_c1,net334_c1);
SPLITT SplitCLK_4_205(net331,net333_c1,net332_c1);
SPLITT SplitCLK_0_206(net298,net330_c1,net331_c1);
SPLITT SplitCLK_0_207(net324,net328_c1,net329_c1);
SPLITT SplitCLK_4_208(net325,net326_c1,net327_c1);
SPLITT SplitCLK_4_209(net316,net324_c1,net325_c1);
SPLITT SplitCLK_0_210(net318,net322_c1,net323_c1);
SPLITT SplitCLK_4_211(net319,net321_c1,net320_c1);
SPLITT SplitCLK_6_212(net317,net318_c1,net319_c1);
SPLITT SplitCLK_6_213(net300,net316_c1,net317_c1);
SPLITT SplitCLK_0_214(net310,net314_c1,net315_c1);
SPLITT SplitCLK_4_215(net311,net312_c1,net313_c1);
SPLITT SplitCLK_0_216(net302,net310_c1,net311_c1);
SPLITT SplitCLK_4_217(net304,net309_c1,net308_c1);
SPLITT SplitCLK_4_218(net305,net307_c1,net306_c1);
SPLITT SplitCLK_6_219(net303,net305_c1,net304_c1);
SPLITT SplitCLK_4_220(net301,net303_c1,net302_c1);
SPLITT SplitCLK_2_221(net299,net301_c1,net300_c1);
SPLITT SplitCLK_6_222(net234,net298_c1,net299_c1);
SPLITT SplitCLK_0_223(net292,net296_c1,net297_c1);
SPLITT SplitCLK_4_224(net293,net294_c1,net295_c1);
SPLITT SplitCLK_0_225(net284,net292_c1,net293_c1);
SPLITT SplitCLK_0_226(net286,net290_c1,net291_c1);
SPLITT SplitCLK_4_227(net287,net288_c1,net289_c1);
SPLITT SplitCLK_6_228(net285,net287_c1,net286_c1);
SPLITT SplitCLK_6_229(net268,net284_c1,net285_c1);
SPLITT SplitCLK_4_230(net278,net282_c1,net283_c1);
SPLITT SplitCLK_4_231(net279,net281_c1,net280_c1);
SPLITT SplitCLK_4_232(net270,net279_c1,net278_c1);
SPLITT SplitCLK_0_233(net272,net277_c1,net276_c1);
SPLITT SplitCLK_4_234(net273,net274_c1,net275_c1);
SPLITT SplitCLK_6_235(net271,net272_c1,net273_c1);
SPLITT SplitCLK_4_236(net269,net271_c1,net270_c1);
SPLITT SplitCLK_4_237(net236,net269_c1,net268_c1);
SPLITT SplitCLK_0_238(net262,net267_c1,net266_c1);
SPLITT SplitCLK_4_239(net263,net265_c1,net264_c1);
SPLITT SplitCLK_0_240(net254,net262_c1,net263_c1);
SPLITT SplitCLK_4_241(net256,net260_c1,net261_c1);
SPLITT SplitCLK_4_242(net257,net258_c1,net259_c1);
SPLITT SplitCLK_6_243(net255,net257_c1,net256_c1);
SPLITT SplitCLK_6_244(net238,net254_c1,net255_c1);
SPLITT SplitCLK_4_245(net248,net253_c1,net252_c1);
SPLITT SplitCLK_4_246(net249,net251_c1,net250_c1);
SPLITT SplitCLK_4_247(net240,net248_c1,net249_c1);
SPLITT SplitCLK_0_248(net242,net246_c1,net247_c1);
SPLITT SplitCLK_4_249(net243,net244_c1,net245_c1);
SPLITT SplitCLK_6_250(net241,net243_c1,net242_c1);
SPLITT SplitCLK_4_251(net239,net241_c1,net240_c1);
SPLITT SplitCLK_2_252(net237,net239_c1,net238_c1);
SPLITT SplitCLK_4_253(net235,net237_c1,net236_c1);
SPLITT SplitCLK_2_254(net233,net235_c1,net234_c1);
SPLITT SplitCLK_0_255(net486,net232_c1,net233_c1);
INTERCONNECT TMS_Pad_Split_136_n349(TMS_Pad,net0);
INTERCONNECT AND2T_16_n40_AND2T_17_n41(net1_c1,net1);
INTERCONNECT NOTT_8_n32_AND2T_63_n93(net2_c1,net2);
INTERCONNECT AND2T_17_n41_Split_146_n359(net3_c1,net3);
INTERCONNECT AND2T_9_n33_DFFT_65__PIPL_n95(net4_c1,net4);
INTERCONNECT OR2T_26_n50_OR2T_27_n51(net5_c1,net5);
INTERCONNECT NOTT_18_n42_Split_147_n360(net6_c1,net6);
INTERCONNECT AND2T_10_n34_DFFT_66__PIPL_n96(net7_c1,net7);
INTERCONNECT OR2T_27_n51_OR2T_34_n58(net8_c1,net8);
INTERCONNECT AND2T_19_n43_Split_148_n361(net9_c1,net9);
INTERCONNECT AND2T_11_n35_Split_139_n352(net10_c1,net10);
INTERCONNECT OR2T_36_n60_Split_162_n375(net11_c1,net11);
INTERCONNECT AND2T_28_n52_Split_156_n369(net12_c1,net12);
INTERCONNECT AND2T_20_n44_Split_149_n362(net13_c1,net13);
INTERCONNECT NOTT_12_n36_Split_140_n353(net14_c1,net14);
INTERCONNECT OR2T_37_n61_AND2T_43_n67(net15_c1,net15);
INTERCONNECT XOR2T_29_n53_DFFT_83__FPB_n296(net16_c1,net16);
INTERCONNECT AND2T_21_n45_OR2T_23_n47(net17_c1,net17);
INTERCONNECT NOTT_13_n37_Split_143_n356(net18_c1,net18);
INTERCONNECT AND2T_46_n70_DFFT_100__FPB_n313(net19_c1,net19);
INTERCONNECT NOTT_38_n62_Split_163_n376(net20_c1,net20);
INTERCONNECT AND2T_30_n54_AND2T_31_n55(net21_c1,net21);
INTERCONNECT AND2T_22_n46_OR2T_23_n47(net22_c1,net22);
INTERCONNECT AND2T_14_n38_Split_144_n357(net23_c1,net23);
INTERCONNECT AND2T_47_n71_OR2T_48_n72(net24_c1,net24);
INTERCONNECT AND2T_39_n63_AND2T_40_n64(net25_c1,net25);
INTERCONNECT AND2T_31_n55_OR2T_32_n56(net26_c1,net26);
INTERCONNECT OR2T_23_n47_Split_151_n364(net27_c1,net27);
INTERCONNECT NOTT_15_n39_Split_145_n358(net28_c1,net28);
INTERCONNECT OR2T_56_n80_DFFT_107__FPB_n320(net29_c1,net29);
INTERCONNECT OR2T_48_n72_AND2T_51_n75(net30_c1,net30);
INTERCONNECT AND2T_40_n64_OR2T_41_n65(net31_c1,net31);
INTERCONNECT OR2T_32_n56_Split_157_n370(net32_c1,net32);
INTERCONNECT AND2T_24_n48_Split_153_n366(net33_c1,net33);
INTERCONNECT AND2T_57_n81_DFFT_71__FBL_n284(net34_c1,net34);
INTERCONNECT OR2T_49_n73_DFFT_101__FPB_n314(net35_c1,net35);
INTERCONNECT OR2T_41_n65_Split_165_n378(net36_c1,net36);
INTERCONNECT OR2T_33_n57_OR2T_34_n58(net37_c1,net37);
INTERCONNECT AND2T_25_n49_Split_154_n367(net38_c1,net38);
INTERCONNECT NOTT_58_n82_DFFT_109__FPB_n322(net39_c1,net39);
INTERCONNECT AND2T_50_n74_AND2T_51_n75(net40_c1,net40);
INTERCONNECT OR2T_42_n66_AND2T_43_n67(net41_c1,net41);
INTERCONNECT OR2T_34_n58_Split_159_n372(net42_c1,net42);
INTERCONNECT AND2T_59_n83_AND2T_60_n84(net43_c1,net43);
INTERCONNECT AND2T_51_n75_OR2T_52_n76(net44_c1,net44);
INTERCONNECT AND2T_43_n67_DFFT_97__FPB_n310(net45_c1,net45);
INTERCONNECT AND2T_35_n59_Split_160_n373(net46_c1,net46);
INTERCONNECT AND2T_60_n84_AND2T_61_n85(net47_c1,net47);
INTERCONNECT OR2T_52_n76_AND2T_53_n77(net48_c1,net48);
INTERCONNECT AND2T_44_n68_Split_166_n379(net49_c1,net49);
INTERCONNECT AND2T_63_n93_Split_169_n382(net50_c1,net50);
INTERCONNECT AND2T_61_n85_DFFT_110__FPB_n323(net51_c1,net51);
INTERCONNECT AND2T_53_n77_Split_168_n381(net52_c1,net52);
INTERCONNECT AND2T_45_n69_Split_167_n380(net53_c1,net53);
INTERCONNECT NOTT_64_n94_Split_172_n385(net54_c1,net54);
INTERCONNECT AND2T_62_n86_DFFT_75__FPB_n288(net55_c1,net55);
INTERCONNECT AND2T_54_n78_OR2T_55_n79(net56_c1,net56);
INTERCONNECT OR2T_55_n79_OR2T_56_n80(net57_c1,net57);
INTERCONNECT Split_137_n350_OR2T_49_n73(net58_c1,net58);
INTERCONNECT Split_138_n351_DFFT_108__FPB_n321(net59_c1,net59);
INTERCONNECT Split_147_n360_DFFT_86__FPB_n299(net60_c1,net60);
INTERCONNECT Split_139_n352_AND2T_60_n84(net61_c1,net61);
INTERCONNECT Split_140_n353_Split_142_n355(net62_c1,net62);
INTERCONNECT Split_148_n361_DFFT_81__FPB_n294(net63_c1,net63);
INTERCONNECT Split_157_n370_Split_158_n371(net64_c1,net64);
INTERCONNECT Split_149_n362_Split_150_n363(net65_c1,net65);
INTERCONNECT Split_141_n354_AND2T_39_n63(net66_c1,net66);
INTERCONNECT Split_142_n355_DFFT_82__FPB_n295(net67_c1,net67);
INTERCONNECT Split_158_n371_OR2T_37_n61(net68_c1,net68);
INTERCONNECT Split_150_n363_AND2T_25_n49(net69_c1,net69);
INTERCONNECT Split_167_n380_DFFT_104__FPB_n317(net70_c1,net70);
INTERCONNECT Split_151_n364_Split_152_n365(net71_c1,net71);
INTERCONNECT Split_159_n372_AND2T_62_n86(net72_c1,net72);
INTERCONNECT Split_143_n356_AND2T_30_n54(net73_c1,net73);
INTERCONNECT Split_136_n349_Split_138_n351(net74_c1,net74);
INTERCONNECT Split_168_n381_DFFT_74__FBL_n287(net75_c1,net75);
INTERCONNECT Split_160_n373_Split_161_n374(net76_c1,net76);
INTERCONNECT Split_152_n365_OR2T_42_n66(net77_c1,net77);
INTERCONNECT Split_144_n357_AND2T_22_n46(net78_c1,net78);
INTERCONNECT Split_169_n382_Split_171_n384(net79_c1,net79);
INTERCONNECT Split_177_n390_Split_178_n391(net80_c1,net80);
INTERCONNECT Split_161_n374_AND2T_53_n77(net81_c1,net81);
INTERCONNECT Split_153_n366_AND2T_54_n78(net82_c1,net82);
INTERCONNECT Split_145_n358_AND2T_20_n44(net83_c1,net83);
INTERCONNECT Split_154_n367_Split_155_n368(net84_c1,net84);
INTERCONNECT Split_162_n375_AND2T_50_n74(net85_c1,net85);
INTERCONNECT Split_146_n359_DFFT_68__PIPL_n98(net86_c1,net86);
INTERCONNECT Split_170_n383_AND2T_24_n48(net87_c1,net87);
INTERCONNECT Split_178_n391_DFFT_78__FPB_n291(net88_c1,net88);
INTERCONNECT Split_163_n376_Split_164_n377(net89_c1,net89);
INTERCONNECT Split_179_n392_Split_180_n393(net90_c1,net90);
INTERCONNECT Split_171_n384_DFFT_67__PIPL_n97(net91_c1,net91);
INTERCONNECT Split_155_n368_OR2T_36_n60(net92_c1,net92);
INTERCONNECT Split_172_n385_Split_174_n387(net93_c1,net93);
INTERCONNECT Split_156_n369_DFFT_98__FPB_n311(net94_c1,net94);
INTERCONNECT Split_164_n377_DFFT_95__FPB_n308(net95_c1,net95);
INTERCONNECT Split_180_n393_NOTT_64_n94(net96_c1,net96);
INTERCONNECT Split_181_n394_Split_183_n396(net97_c1,net97);
INTERCONNECT Split_165_n378_AND2T_45_n69(net98_c1,net98);
INTERCONNECT Split_173_n386_AND2T_10_n34(net99_c1,net99);
INTERCONNECT TRST_Pad_NOTT_18_n42(TRST_Pad,net100);
INTERCONNECT Split_166_n379_DFFT_73__FBL_n286(net101_c1,net101);
INTERCONNECT Split_182_n395_AND2T_19_n43(net102_c1,net102);
INTERCONNECT Split_174_n387_AND2T_20_n44(net103_c1,net103);
INTERCONNECT Split_175_n388_Split_176_n389(net104_c1,net104);
INTERCONNECT Split_183_n396_DFFT_76__FPB_n289(net105_c1,net105);
INTERCONNECT Split_184_n397_Split_186_n399(net106_c1,net106);
INTERCONNECT Split_176_n389_DFFT_94__FPB_n307(net107_c1,net107);
INTERCONNECT Split_185_n398_AND2T_19_n43(net108_c1,net108);
INTERCONNECT Split_186_n399_DFFT_77__FPB_n290(net109_c1,net109);
INTERCONNECT Split_137_n350_NOTT_38_n62(net110_c1,net110);
INTERCONNECT Split_138_n351_DFFT_91__FPB_n304(net111_c1,net111);
INTERCONNECT Split_139_n352_AND2T_40_n64(net112_c1,net112);
INTERCONNECT Split_147_n360_AND2T_59_n83(net113_c1,net113);
INTERCONNECT Split_148_n361_DFFT_80__FPB_n293(net114_c1,net114);
INTERCONNECT Split_140_n353_Split_141_n354(net115_c1,net115);
INTERCONNECT Split_149_n362_AND2T_31_n55(net116_c1,net116);
INTERCONNECT Split_157_n370_OR2T_48_n72(net117_c1,net117);
INTERCONNECT Split_141_n354_AND2T_14_n38(net118_c1,net118);
INTERCONNECT Split_158_n371_OR2T_33_n57(net119_c1,net119);
INTERCONNECT Split_142_n355_NOTT_58_n82(net120_c1,net120);
INTERCONNECT Split_150_n363_AND2T_21_n45(net121_c1,net121);
INTERCONNECT Split_159_n372_AND2T_35_n59(net122_c1,net122);
INTERCONNECT Split_167_n380_OR2T_56_n80(net123_c1,net123);
INTERCONNECT Split_143_n356_AND2T_14_n38(net124_c1,net124);
INTERCONNECT Split_151_n364_OR2T_55_n79(net125_c1,net125);
INTERCONNECT Split_168_n381_DFFT_70__FBL_n283(net126_c1,net126);
INTERCONNECT Split_136_n349_Split_137_n350(net127_c1,net127);
INTERCONNECT Split_144_n357_AND2T_17_n41(net128_c1,net128);
INTERCONNECT Split_152_n365_OR2T_27_n51(net129_c1,net129);
INTERCONNECT Split_160_n373_AND2T_57_n81(net130_c1,net130);
INTERCONNECT Split_169_n382_Split_170_n383(net131_c1,net131);
INTERCONNECT Split_177_n390_DFFT_112__FPB_n325(net132_c1,net132);
INTERCONNECT Split_145_n358_AND2T_16_n40(net133_c1,net133);
INTERCONNECT Split_153_n366_OR2T_26_n50(net134_c1,net134);
INTERCONNECT Split_161_n374_AND2T_44_n68(net135_c1,net135);
INTERCONNECT Split_178_n391_NOTT_15_n39(net136_c1,net136);
INTERCONNECT Split_146_n359_OR2T_32_n56(net137_c1,net137);
INTERCONNECT Split_154_n367_AND2T_47_n71(net138_c1,net138);
INTERCONNECT Split_162_n375_OR2T_37_n61(net139_c1,net139);
INTERCONNECT Split_170_n383_AND2T_22_n46(net140_c1,net140);
INTERCONNECT Split_179_n392_DFFT_79__FPB_n292(net141_c1,net141);
INTERCONNECT Split_155_n368_OR2T_26_n50(net142_c1,net142);
INTERCONNECT Split_163_n376_DFFT_105__FPB_n318(net143_c1,net143);
INTERCONNECT Split_171_n384_AND2T_28_n52(net144_c1,net144);
INTERCONNECT Split_156_n369_DFFT_85__FPB_n298(net145_c1,net145);
INTERCONNECT Split_164_n377_AND2T_46_n70(net146_c1,net146);
INTERCONNECT Split_172_n385_Split_173_n386(net147_c1,net147);
INTERCONNECT Split_180_n393_NOTT_8_n32(net148_c1,net148);
INTERCONNECT Split_165_n378_OR2T_42_n66(net149_c1,net149);
INTERCONNECT Split_173_n386_AND2T_9_n33(net150_c1,net150);
INTERCONNECT Split_181_n394_Split_182_n395(net151_c1,net151);
INTERCONNECT Split_166_n379_DFFT_69__FBL_n282(net152_c1,net152);
INTERCONNECT Split_174_n387_AND2T_11_n35(net153_c1,net153);
INTERCONNECT Split_182_n395_NOTT_12_n36(net154_c1,net154);
INTERCONNECT Split_175_n388_DFFT_99__FPB_n312(net155_c1,net155);
INTERCONNECT Split_183_n396_XOR2T_29_n53(net156_c1,net156);
INTERCONNECT Split_176_n389_OR2T_49_n73(net157_c1,net157);
INTERCONNECT Split_184_n397_Split_185_n398(net158_c1,net158);
INTERCONNECT Split_185_n398_NOTT_13_n37(net159_c1,net159);
INTERCONNECT Split_186_n399_XOR2T_29_n53(net160_c1,net160);
INTERCONNECT DFFT_69__FBL_n282_DFFT_84__FPB_n297(net161_c1,net161);
INTERCONNECT DFFT_70__FBL_n283_Split_175_n388(net162_c1,net162);
INTERCONNECT DFFT_71__FBL_n284_Split_177_n390(net163_c1,net163);
INTERCONNECT DFFT_72__FBL_n285_Split_179_n392(net164_c1,net164);
INTERCONNECT DFFT_73__FBL_n286_Split_181_n394(net165_c1,net165);
INTERCONNECT DFFT_74__FBL_n287_Split_184_n397(net166_c1,net166);
INTERCONNECT DFFT_87__FPB_n300_DFFT_88__FPB_n301(net167_c1,net167);
INTERCONNECT DFFT_88__FPB_n301_DFFT_89__FPB_n302(net168_c1,net168);
INTERCONNECT DFFT_89__FPB_n302_DFFT_90__FPB_n303(net169_c1,net169);
INTERCONNECT DFFT_97__FPB_n310_AND2T_44_n68(net170_c1,net170);
INTERCONNECT DFFT_98__FPB_n311_AND2T_45_n69(net171_c1,net171);
INTERCONNECT DFFT_90__FPB_n303_AND2T_35_n59(net172_c1,net172);
INTERCONNECT DFFT_91__FPB_n304_DFFT_92__FPB_n305(net173_c1,net173);
INTERCONNECT DFFT_107__FPB_n320_AND2T_57_n81(net174_c1,net174);
INTERCONNECT DFFT_99__FPB_n312_AND2T_46_n70(net175_c1,net175);
INTERCONNECT DFFT_92__FPB_n305_DFFT_93__FPB_n306(net176_c1,net176);
INTERCONNECT DFFT_108__FPB_n321_AND2T_59_n83(net177_c1,net177);
INTERCONNECT DFFT_100__FPB_n313_AND2T_47_n71(net178_c1,net178);
INTERCONNECT DFFT_117__FPB_n330_DFFT_118_state_obs0(net179_c1,net179);
INTERCONNECT DFFT_101__FPB_n314_DFFT_102__FPB_n315(net180_c1,net180);
INTERCONNECT DFFT_109__FPB_n322_AND2T_61_n85(net181_c1,net181);
INTERCONNECT DFFT_93__FPB_n306_OR2T_36_n60(net182_c1,net182);
INTERCONNECT DFFT_110__FPB_n323_DFFT_111__FPB_n324(net183_c1,net183);
INTERCONNECT DFFT_102__FPB_n315_DFFT_103__FPB_n316(net184_c1,net184);
INTERCONNECT DFFT_94__FPB_n307_AND2T_39_n63(net185_c1,net185);
INTERCONNECT DFFT_127__FPB_n340_DFFT_128__FPB_n341(net186_c1,net186);
INTERCONNECT DFFT_119__FPB_n332_DFFT_120__FPB_n333(net187_c1,net187);
INTERCONNECT DFFT_95__FPB_n308_DFFT_96__FPB_n309(net188_c1,net188);
INTERCONNECT DFFT_111__FPB_n324_AND2T_62_n86(net189_c1,net189);
INTERCONNECT DFFT_103__FPB_n316_AND2T_50_n74(net190_c1,net190);
INTERCONNECT DFFT_128__FPB_n341_DFFT_129__FPB_n342(net191_c1,net191);
INTERCONNECT DFFT_120__FPB_n333_DFFT_121__FPB_n334(net192_c1,net192);
INTERCONNECT DFFT_112__FPB_n325_AND2T_63_n93(net193_c1,net193);
INTERCONNECT DFFT_104__FPB_n317_OR2T_52_n76(net194_c1,net194);
INTERCONNECT DFFT_96__FPB_n309_OR2T_41_n65(net195_c1,net195);
INTERCONNECT DFFT_129__FPB_n342_DFFT_130_state_obs2(net196_c1,net196);
INTERCONNECT DFFT_121__FPB_n334_DFFT_122__FPB_n335(net197_c1,net197);
INTERCONNECT DFFT_113__FPB_n326_DFFT_114__FPB_n327(net198_c1,net198);
INTERCONNECT DFFT_105__FPB_n318_DFFT_106__FPB_n319(net199_c1,net199);
INTERCONNECT DFFT_122__FPB_n335_DFFT_123__FPB_n336(net200_c1,net200);
INTERCONNECT DFFT_114__FPB_n327_DFFT_115__FPB_n328(net201_c1,net201);
INTERCONNECT DFFT_106__FPB_n319_AND2T_54_n78(net202_c1,net202);
INTERCONNECT DFFT_131__FPB_n344_DFFT_132__FPB_n345(net203_c1,net203);
INTERCONNECT DFFT_123__FPB_n336_DFFT_124_state_obs1(net204_c1,net204);
INTERCONNECT DFFT_115__FPB_n328_DFFT_116__FPB_n329(net205_c1,net205);
INTERCONNECT DFFT_132__FPB_n345_DFFT_133__FPB_n346(net206_c1,net206);
INTERCONNECT DFFT_116__FPB_n329_DFFT_117__FPB_n330(net207_c1,net207);
INTERCONNECT DFFT_133__FPB_n346_DFFT_134__FPB_n347(net208_c1,net208);
INTERCONNECT DFFT_125__FPB_n338_DFFT_126__FPB_n339(net209_c1,net209);
INTERCONNECT DFFT_77__FPB_n290_AND2T_10_n34(net210_c1,net210);
INTERCONNECT DFFT_134__FPB_n347_DFFT_135_state_obs3(net211_c1,net211);
INTERCONNECT DFFT_126__FPB_n339_DFFT_127__FPB_n340(net212_c1,net212);
INTERCONNECT DFFT_78__FPB_n291_AND2T_11_n35(net213_c1,net213);
INTERCONNECT DFFT_79__FPB_n292_AND2T_16_n40(net214_c1,net214);
INTERCONNECT DFFT_80__FPB_n293_AND2T_21_n45(net215_c1,net215);
INTERCONNECT DFFT_81__FPB_n294_AND2T_24_n48(net216_c1,net216);
INTERCONNECT DFFT_82__FPB_n295_AND2T_25_n49(net217_c1,net217);
INTERCONNECT DFFT_75__FPB_n288_DFFT_72__FBL_n285(net218_c1,net218);
INTERCONNECT DFFT_83__FPB_n296_AND2T_28_n52(net219_c1,net219);
INTERCONNECT DFFT_84__FPB_n297_AND2T_30_n54(net220_c1,net220);
INTERCONNECT DFFT_76__FPB_n289_AND2T_9_n33(net221_c1,net221);
INTERCONNECT DFFT_85__FPB_n298_OR2T_33_n57(net222_c1,net222);
INTERCONNECT DFFT_86__FPB_n299_DFFT_87__FPB_n300(net223_c1,net223);
INTERCONNECT DFFT_65__PIPL_n95_DFFT_113__FPB_n326(net224_c1,net224);
INTERCONNECT DFFT_66__PIPL_n96_DFFT_119__FPB_n332(net225_c1,net225);
INTERCONNECT DFFT_67__PIPL_n97_DFFT_125__FPB_n338(net226_c1,net226);
INTERCONNECT DFFT_68__PIPL_n98_DFFT_131__FPB_n344(net227_c1,net227);
INTERCONNECT DFFT_118_state_obs0_state_obs0_Pad(net228_c1,state_obs0_Pad);
INTERCONNECT DFFT_124_state_obs1_state_obs1_Pad(net229_c1,state_obs1_Pad);
INTERCONNECT DFFT_130_state_obs2_state_obs2_Pad(net230_c1,state_obs2_Pad);
INTERCONNECT DFFT_135_state_obs3_state_obs3_Pad(net231_c1,state_obs3_Pad);
INTERCONNECT SplitCLK_0_255_SplitCLK_0_191(net232_c1,net232);
INTERCONNECT SplitCLK_0_255_SplitCLK_2_254(net233_c1,net233);
INTERCONNECT SplitCLK_2_254_SplitCLK_6_222(net234_c1,net234);
INTERCONNECT SplitCLK_2_254_SplitCLK_4_253(net235_c1,net235);
INTERCONNECT SplitCLK_4_253_SplitCLK_4_237(net236_c1,net236);
INTERCONNECT SplitCLK_4_253_SplitCLK_2_252(net237_c1,net237);
INTERCONNECT SplitCLK_2_252_SplitCLK_6_244(net238_c1,net238);
INTERCONNECT SplitCLK_2_252_SplitCLK_4_251(net239_c1,net239);
INTERCONNECT SplitCLK_4_251_SplitCLK_4_247(net240_c1,net240);
INTERCONNECT SplitCLK_4_251_SplitCLK_6_250(net241_c1,net241);
INTERCONNECT SplitCLK_6_250_SplitCLK_0_248(net242_c1,net242);
INTERCONNECT SplitCLK_6_250_SplitCLK_4_249(net243_c1,net243);
INTERCONNECT SplitCLK_4_249_OR2T_49_n73(net244_c1,net244);
INTERCONNECT SplitCLK_4_249_DFFT_101__FPB_n314(net245_c1,net245);
INTERCONNECT SplitCLK_0_248_OR2T_52_n76(net246_c1,net246);
INTERCONNECT SplitCLK_0_248_DFFT_70__FBL_n283(net247_c1,net247);
INTERCONNECT SplitCLK_4_247_SplitCLK_4_245(net248_c1,net248);
INTERCONNECT SplitCLK_4_247_SplitCLK_4_246(net249_c1,net249);
INTERCONNECT SplitCLK_4_246_DFFT_102__FPB_n315(net250_c1,net250);
INTERCONNECT SplitCLK_4_246_DFFT_108__FPB_n321(net251_c1,net251);
INTERCONNECT SplitCLK_4_245_DFFT_103__FPB_n316(net252_c1,net252);
INTERCONNECT SplitCLK_4_245_DFFT_104__FPB_n317(net253_c1,net253);
INTERCONNECT SplitCLK_6_244_SplitCLK_0_240(net254_c1,net254);
INTERCONNECT SplitCLK_6_244_SplitCLK_6_243(net255_c1,net255);
INTERCONNECT SplitCLK_6_243_SplitCLK_4_241(net256_c1,net256);
INTERCONNECT SplitCLK_6_243_SplitCLK_4_242(net257_c1,net257);
INTERCONNECT SplitCLK_4_242_AND2T_44_n68(net258_c1,net258);
INTERCONNECT SplitCLK_4_242_AND2T_53_n77(net259_c1,net259);
INTERCONNECT SplitCLK_4_241_NOTT_12_n36(net260_c1,net260);
INTERCONNECT SplitCLK_4_241_DFFT_97__FPB_n310(net261_c1,net261);
INTERCONNECT SplitCLK_0_240_SplitCLK_0_238(net262_c1,net262);
INTERCONNECT SplitCLK_0_240_SplitCLK_4_239(net263_c1,net263);
INTERCONNECT SplitCLK_4_239_AND2T_51_n75(net264_c1,net264);
INTERCONNECT SplitCLK_4_239_AND2T_43_n67(net265_c1,net265);
INTERCONNECT SplitCLK_0_238_OR2T_33_n57(net266_c1,net266);
INTERCONNECT SplitCLK_0_238_DFFT_74__FBL_n287(net267_c1,net267);
INTERCONNECT SplitCLK_4_237_SplitCLK_6_229(net268_c1,net268);
INTERCONNECT SplitCLK_4_237_SplitCLK_4_236(net269_c1,net269);
INTERCONNECT SplitCLK_4_236_SplitCLK_4_232(net270_c1,net270);
INTERCONNECT SplitCLK_4_236_SplitCLK_6_235(net271_c1,net271);
INTERCONNECT SplitCLK_6_235_SplitCLK_0_233(net272_c1,net272);
INTERCONNECT SplitCLK_6_235_SplitCLK_4_234(net273_c1,net273);
INTERCONNECT SplitCLK_4_234_DFFT_91__FPB_n304(net274_c1,net274);
INTERCONNECT SplitCLK_4_234_DFFT_92__FPB_n305(net275_c1,net275);
INTERCONNECT SplitCLK_0_233_AND2T_50_n74(net276_c1,net276);
INTERCONNECT SplitCLK_0_233_OR2T_37_n61(net277_c1,net277);
INTERCONNECT SplitCLK_4_232_SplitCLK_4_230(net278_c1,net278);
INTERCONNECT SplitCLK_4_232_SplitCLK_4_231(net279_c1,net279);
INTERCONNECT SplitCLK_4_231_NOTT_38_n62(net280_c1,net280);
INTERCONNECT SplitCLK_4_231_DFFT_93__FPB_n306(net281_c1,net281);
INTERCONNECT SplitCLK_4_230_DFFT_94__FPB_n307(net282_c1,net282);
INTERCONNECT SplitCLK_4_230_DFFT_89__FPB_n302(net283_c1,net283);
INTERCONNECT SplitCLK_6_229_SplitCLK_0_225(net284_c1,net284);
INTERCONNECT SplitCLK_6_229_SplitCLK_6_228(net285_c1,net285);
INTERCONNECT SplitCLK_6_228_SplitCLK_0_226(net286_c1,net286);
INTERCONNECT SplitCLK_6_228_SplitCLK_4_227(net287_c1,net287);
INTERCONNECT SplitCLK_4_227_AND2T_45_n69(net288_c1,net288);
INTERCONNECT SplitCLK_4_227_AND2T_39_n63(net289_c1,net289);
INTERCONNECT SplitCLK_0_226_DFFT_85__FPB_n298(net290_c1,net290);
INTERCONNECT SplitCLK_0_226_DFFT_98__FPB_n311(net291_c1,net291);
INTERCONNECT SplitCLK_0_225_SplitCLK_0_223(net292_c1,net292);
INTERCONNECT SplitCLK_0_225_SplitCLK_4_224(net293_c1,net293);
INTERCONNECT SplitCLK_4_224_OR2T_42_n66(net294_c1,net294);
INTERCONNECT SplitCLK_4_224_OR2T_48_n72(net295_c1,net295);
INTERCONNECT SplitCLK_0_223_AND2T_21_n45(net296_c1,net296);
INTERCONNECT SplitCLK_0_223_DFFT_107__FPB_n320(net297_c1,net297);
INTERCONNECT SplitCLK_6_222_SplitCLK_0_206(net298_c1,net298);
INTERCONNECT SplitCLK_6_222_SplitCLK_2_221(net299_c1,net299);
INTERCONNECT SplitCLK_2_221_SplitCLK_6_213(net300_c1,net300);
INTERCONNECT SplitCLK_2_221_SplitCLK_4_220(net301_c1,net301);
INTERCONNECT SplitCLK_4_220_SplitCLK_0_216(net302_c1,net302);
INTERCONNECT SplitCLK_4_220_SplitCLK_6_219(net303_c1,net303);
INTERCONNECT SplitCLK_6_219_SplitCLK_4_217(net304_c1,net304);
INTERCONNECT SplitCLK_6_219_SplitCLK_4_218(net305_c1,net305);
INTERCONNECT SplitCLK_4_218_AND2T_19_n43(net306_c1,net306);
INTERCONNECT SplitCLK_4_218_DFFT_73__FBL_n286(net307_c1,net307);
INTERCONNECT SplitCLK_4_217_NOTT_15_n39(net308_c1,net308);
INTERCONNECT SplitCLK_4_217_DFFT_76__FPB_n289(net309_c1,net309);
INTERCONNECT SplitCLK_0_216_SplitCLK_0_214(net310_c1,net310);
INTERCONNECT SplitCLK_0_216_SplitCLK_4_215(net311_c1,net311);
INTERCONNECT SplitCLK_4_215_AND2T_14_n38(net312_c1,net312);
INTERCONNECT SplitCLK_4_215_AND2T_16_n40(net313_c1,net313);
INTERCONNECT SplitCLK_0_214_AND2T_9_n33(net314_c1,net314);
INTERCONNECT SplitCLK_0_214_AND2T_10_n34(net315_c1,net315);
INTERCONNECT SplitCLK_6_213_SplitCLK_4_209(net316_c1,net316);
INTERCONNECT SplitCLK_6_213_SplitCLK_6_212(net317_c1,net317);
INTERCONNECT SplitCLK_6_212_SplitCLK_0_210(net318_c1,net318);
INTERCONNECT SplitCLK_6_212_SplitCLK_4_211(net319_c1,net319);
INTERCONNECT SplitCLK_4_211_DFFT_114__FPB_n327(net320_c1,net320);
INTERCONNECT SplitCLK_4_211_DFFT_115__FPB_n328(net321_c1,net321);
INTERCONNECT SplitCLK_0_210_DFFT_117__FPB_n330(net322_c1,net322);
INTERCONNECT SplitCLK_0_210_DFFT_118_state_obs0(net323_c1,net323);
INTERCONNECT SplitCLK_4_209_SplitCLK_0_207(net324_c1,net324);
INTERCONNECT SplitCLK_4_209_SplitCLK_4_208(net325_c1,net325);
INTERCONNECT SplitCLK_4_208_DFFT_113__FPB_n326(net326_c1,net326);
INTERCONNECT SplitCLK_4_208_DFFT_65__PIPL_n95(net327_c1,net327);
INTERCONNECT SplitCLK_0_207_DFFT_116__FPB_n329(net328_c1,net328);
INTERCONNECT SplitCLK_0_207_DFFT_124_state_obs1(net329_c1,net329);
INTERCONNECT SplitCLK_0_206_SplitCLK_6_198(net330_c1,net330);
INTERCONNECT SplitCLK_0_206_SplitCLK_4_205(net331_c1,net331);
INTERCONNECT SplitCLK_4_205_SplitCLK_0_201(net332_c1,net332);
INTERCONNECT SplitCLK_4_205_SplitCLK_2_204(net333_c1,net333);
INTERCONNECT SplitCLK_2_204_SplitCLK_4_202(net334_c1,net334);
INTERCONNECT SplitCLK_2_204_SplitCLK_4_203(net335_c1,net335);
INTERCONNECT SplitCLK_4_203_NOTT_13_n37(net336_c1,net336);
INTERCONNECT SplitCLK_4_203_DFFT_81__FPB_n294(net337_c1,net337);
INTERCONNECT SplitCLK_4_202_AND2T_20_n44(net338_c1,net338);
INTERCONNECT SplitCLK_4_202_DFFT_77__FPB_n290(net339_c1,net339);
INTERCONNECT SplitCLK_0_201_SplitCLK_4_199(net340_c1,net340);
INTERCONNECT SplitCLK_0_201_SplitCLK_4_200(net341_c1,net341);
INTERCONNECT SplitCLK_4_200_DFFT_80__FPB_n293(net342_c1,net342);
INTERCONNECT SplitCLK_4_200_DFFT_69__FBL_n282(net343_c1,net343);
INTERCONNECT SplitCLK_4_199_XOR2T_29_n53(net344_c1,net344);
INTERCONNECT SplitCLK_4_199_AND2T_17_n41(net345_c1,net345);
INTERCONNECT SplitCLK_6_198_SplitCLK_4_194(net346_c1,net346);
INTERCONNECT SplitCLK_6_198_SplitCLK_6_197(net347_c1,net347);
INTERCONNECT SplitCLK_6_197_SplitCLK_0_195(net348_c1,net348);
INTERCONNECT SplitCLK_6_197_SplitCLK_4_196(net349_c1,net349);
INTERCONNECT SplitCLK_4_196_DFFT_119__FPB_n332(net350_c1,net350);
INTERCONNECT SplitCLK_4_196_DFFT_66__PIPL_n96(net351_c1,net351);
INTERCONNECT SplitCLK_0_195_DFFT_122__FPB_n335(net352_c1,net352);
INTERCONNECT SplitCLK_0_195_DFFT_123__FPB_n336(net353_c1,net353);
INTERCONNECT SplitCLK_4_194_SplitCLK_0_192(net354_c1,net354);
INTERCONNECT SplitCLK_4_194_SplitCLK_4_193(net355_c1,net355);
INTERCONNECT SplitCLK_4_193_DFFT_120__FPB_n333(net356_c1,net356);
INTERCONNECT SplitCLK_4_193_DFFT_121__FPB_n334(net357_c1,net357);
INTERCONNECT SplitCLK_0_192_DFFT_129__FPB_n342(net358_c1,net358);
INTERCONNECT SplitCLK_0_192_DFFT_130_state_obs2(net359_c1,net359);
INTERCONNECT SplitCLK_0_191_SplitCLK_6_159(net360_c1,net360);
INTERCONNECT SplitCLK_0_191_SplitCLK_4_190(net361_c1,net361);
INTERCONNECT SplitCLK_4_190_SplitCLK_0_174(net362_c1,net362);
INTERCONNECT SplitCLK_4_190_SplitCLK_2_189(net363_c1,net363);
INTERCONNECT SplitCLK_2_189_SplitCLK_2_181(net364_c1,net364);
INTERCONNECT SplitCLK_2_189_SplitCLK_4_188(net365_c1,net365);
INTERCONNECT SplitCLK_4_188_SplitCLK_0_184(net366_c1,net366);
INTERCONNECT SplitCLK_4_188_SplitCLK_2_187(net367_c1,net367);
INTERCONNECT SplitCLK_2_187_SplitCLK_4_185(net368_c1,net368);
INTERCONNECT SplitCLK_2_187_SplitCLK_4_186(net369_c1,net369);
INTERCONNECT SplitCLK_4_186_DFFT_90__FPB_n303(net370_c1,net370);
INTERCONNECT SplitCLK_4_186_DFFT_88__FPB_n301(net371_c1,net371);
INTERCONNECT SplitCLK_4_185_DFFT_99__FPB_n312(net372_c1,net372);
INTERCONNECT SplitCLK_4_185_OR2T_36_n60(net373_c1,net373);
INTERCONNECT SplitCLK_0_184_SplitCLK_0_182(net374_c1,net374);
INTERCONNECT SplitCLK_0_184_SplitCLK_4_183(net375_c1,net375);
INTERCONNECT SplitCLK_4_183_DFFT_86__FPB_n299(net376_c1,net376);
INTERCONNECT SplitCLK_4_183_DFFT_87__FPB_n300(net377_c1,net377);
INTERCONNECT SplitCLK_0_182_AND2T_46_n70(net378_c1,net378);
INTERCONNECT SplitCLK_0_182_DFFT_100__FPB_n313(net379_c1,net379);
INTERCONNECT SplitCLK_2_181_SplitCLK_4_177(net380_c1,net380);
INTERCONNECT SplitCLK_2_181_SplitCLK_2_180(net381_c1,net381);
INTERCONNECT SplitCLK_2_180_SplitCLK_4_178(net382_c1,net382);
INTERCONNECT SplitCLK_2_180_SplitCLK_4_179(net383_c1,net383);
INTERCONNECT SplitCLK_4_179_AND2T_47_n71(net384_c1,net384);
INTERCONNECT SplitCLK_4_179_OR2T_56_n80(net385_c1,net385);
INTERCONNECT SplitCLK_4_178_AND2T_57_n81(net386_c1,net386);
INTERCONNECT SplitCLK_4_178_OR2T_23_n47(net387_c1,net387);
INTERCONNECT SplitCLK_4_177_SplitCLK_4_175(net388_c1,net388);
INTERCONNECT SplitCLK_4_177_SplitCLK_4_176(net389_c1,net389);
INTERCONNECT SplitCLK_4_176_AND2T_35_n59(net390_c1,net390);
INTERCONNECT SplitCLK_4_176_OR2T_55_n79(net391_c1,net391);
INTERCONNECT SplitCLK_4_175_OR2T_34_n58(net392_c1,net392);
INTERCONNECT SplitCLK_4_175_DFFT_109__FPB_n322(net393_c1,net393);
INTERCONNECT SplitCLK_0_174_SplitCLK_0_166(net394_c1,net394);
INTERCONNECT SplitCLK_0_174_SplitCLK_4_173(net395_c1,net395);
INTERCONNECT SplitCLK_4_173_SplitCLK_0_169(net396_c1,net396);
INTERCONNECT SplitCLK_4_173_SplitCLK_2_172(net397_c1,net397);
INTERCONNECT SplitCLK_2_172_SplitCLK_4_170(net398_c1,net398);
INTERCONNECT SplitCLK_2_172_SplitCLK_4_171(net399_c1,net399);
INTERCONNECT SplitCLK_4_171_NOTT_18_n42(net400_c1,net400);
INTERCONNECT SplitCLK_4_171_DFFT_106__FPB_n319(net401_c1,net401);
INTERCONNECT SplitCLK_4_170_OR2T_26_n50(net402_c1,net402);
INTERCONNECT SplitCLK_4_170_DFFT_105__FPB_n318(net403_c1,net403);
INTERCONNECT SplitCLK_0_169_SplitCLK_0_167(net404_c1,net404);
INTERCONNECT SplitCLK_0_169_SplitCLK_4_168(net405_c1,net405);
INTERCONNECT SplitCLK_4_168_AND2T_59_n83(net406_c1,net406);
INTERCONNECT SplitCLK_4_168_DFFT_95__FPB_n308(net407_c1,net407);
INTERCONNECT SplitCLK_0_167_AND2T_40_n64(net408_c1,net408);
INTERCONNECT SplitCLK_0_167_AND2T_54_n78(net409_c1,net409);
INTERCONNECT SplitCLK_0_166_SplitCLK_4_162(net410_c1,net410);
INTERCONNECT SplitCLK_0_166_SplitCLK_6_165(net411_c1,net411);
INTERCONNECT SplitCLK_6_165_SplitCLK_4_163(net412_c1,net412);
INTERCONNECT SplitCLK_6_165_SplitCLK_4_164(net413_c1,net413);
INTERCONNECT SplitCLK_4_164_AND2T_61_n85(net414_c1,net414);
INTERCONNECT SplitCLK_4_164_OR2T_27_n51(net415_c1,net415);
INTERCONNECT SplitCLK_4_163_DFFT_110__FPB_n323(net416_c1,net416);
INTERCONNECT SplitCLK_4_163_DFFT_111__FPB_n324(net417_c1,net417);
INTERCONNECT SplitCLK_4_162_SplitCLK_4_160(net418_c1,net418);
INTERCONNECT SplitCLK_4_162_SplitCLK_4_161(net419_c1,net419);
INTERCONNECT SplitCLK_4_161_OR2T_41_n65(net420_c1,net420);
INTERCONNECT SplitCLK_4_161_DFFT_96__FPB_n309(net421_c1,net421);
INTERCONNECT SplitCLK_4_160_AND2T_60_n84(net422_c1,net422);
INTERCONNECT SplitCLK_4_160_AND2T_62_n86(net423_c1,net423);
INTERCONNECT SplitCLK_6_159_SplitCLK_0_143(net424_c1,net424);
INTERCONNECT SplitCLK_6_159_SplitCLK_6_158(net425_c1,net425);
INTERCONNECT SplitCLK_6_158_SplitCLK_6_150(net426_c1,net426);
INTERCONNECT SplitCLK_6_158_SplitCLK_4_157(net427_c1,net427);
INTERCONNECT SplitCLK_4_157_SplitCLK_4_153(net428_c1,net428);
INTERCONNECT SplitCLK_4_157_SplitCLK_2_156(net429_c1,net429);
INTERCONNECT SplitCLK_2_156_SplitCLK_4_154(net430_c1,net430);
INTERCONNECT SplitCLK_2_156_SplitCLK_4_155(net431_c1,net431);
INTERCONNECT SplitCLK_4_155_AND2T_11_n35(net432_c1,net432);
INTERCONNECT SplitCLK_4_155_OR2T_32_n56(net433_c1,net433);
INTERCONNECT SplitCLK_4_154_DFFT_83__FPB_n296(net434_c1,net434);
INTERCONNECT SplitCLK_4_154_DFFT_78__FPB_n291(net435_c1,net435);
INTERCONNECT SplitCLK_4_153_SplitCLK_0_151(net436_c1,net436);
INTERCONNECT SplitCLK_4_153_SplitCLK_4_152(net437_c1,net437);
INTERCONNECT SplitCLK_4_152_AND2T_24_n48(net438_c1,net438);
INTERCONNECT SplitCLK_4_152_AND2T_25_n49(net439_c1,net439);
INTERCONNECT SplitCLK_0_151_AND2T_30_n54(net440_c1,net440);
INTERCONNECT SplitCLK_0_151_AND2T_31_n55(net441_c1,net441);
INTERCONNECT SplitCLK_6_150_SplitCLK_4_146(net442_c1,net442);
INTERCONNECT SplitCLK_6_150_SplitCLK_6_149(net443_c1,net443);
INTERCONNECT SplitCLK_6_149_SplitCLK_4_147(net444_c1,net444);
INTERCONNECT SplitCLK_6_149_SplitCLK_4_148(net445_c1,net445);
INTERCONNECT SplitCLK_4_148_AND2T_28_n52(net446_c1,net446);
INTERCONNECT SplitCLK_4_148_DFFT_125__FPB_n338(net447_c1,net447);
INTERCONNECT SplitCLK_4_147_DFFT_128__FPB_n341(net448_c1,net448);
INTERCONNECT SplitCLK_4_147_DFFT_67__PIPL_n97(net449_c1,net449);
INTERCONNECT SplitCLK_4_146_SplitCLK_4_144(net450_c1,net450);
INTERCONNECT SplitCLK_4_146_SplitCLK_4_145(net451_c1,net451);
INTERCONNECT SplitCLK_4_145_DFFT_126__FPB_n339(net452_c1,net452);
INTERCONNECT SplitCLK_4_145_DFFT_127__FPB_n340(net453_c1,net453);
INTERCONNECT SplitCLK_4_144_DFFT_68__PIPL_n98(net454_c1,net454);
INTERCONNECT SplitCLK_4_144_DFFT_135_state_obs3(net455_c1,net455);
INTERCONNECT SplitCLK_0_143_SplitCLK_6_135(net456_c1,net456);
INTERCONNECT SplitCLK_0_143_SplitCLK_4_142(net457_c1,net457);
INTERCONNECT SplitCLK_4_142_SplitCLK_4_138(net458_c1,net458);
INTERCONNECT SplitCLK_4_142_SplitCLK_2_141(net459_c1,net459);
INTERCONNECT SplitCLK_2_141_SplitCLK_4_139(net460_c1,net460);
INTERCONNECT SplitCLK_2_141_SplitCLK_4_140(net461_c1,net461);
INTERCONNECT SplitCLK_4_140_DFFT_71__FBL_n284(net462_c1,net462);
INTERCONNECT SplitCLK_4_140_DFFT_82__FPB_n295(net463_c1,net463);
INTERCONNECT SplitCLK_4_139_DFFT_112__FPB_n325(net464_c1,net464);
INTERCONNECT SplitCLK_4_139_DFFT_84__FPB_n297(net465_c1,net465);
INTERCONNECT SplitCLK_4_138_SplitCLK_4_136(net466_c1,net466);
INTERCONNECT SplitCLK_4_138_SplitCLK_4_137(net467_c1,net467);
INTERCONNECT SplitCLK_4_137_NOTT_58_n82(net468_c1,net468);
INTERCONNECT SplitCLK_4_137_DFFT_75__FPB_n288(net469_c1,net469);
INTERCONNECT SplitCLK_4_136_AND2T_22_n46(net470_c1,net470);
INTERCONNECT SplitCLK_4_136_DFFT_79__FPB_n292(net471_c1,net471);
INTERCONNECT SplitCLK_6_135_SplitCLK_4_131(net472_c1,net472);
INTERCONNECT SplitCLK_6_135_SplitCLK_6_134(net473_c1,net473);
INTERCONNECT SplitCLK_6_134_SplitCLK_0_132(net474_c1,net474);
INTERCONNECT SplitCLK_6_134_SplitCLK_4_133(net475_c1,net475);
INTERCONNECT SplitCLK_4_133_NOTT_8_n32(net476_c1,net476);
INTERCONNECT SplitCLK_4_133_AND2T_63_n93(net477_c1,net477);
INTERCONNECT SplitCLK_0_132_DFFT_131__FPB_n344(net478_c1,net478);
INTERCONNECT SplitCLK_0_132_DFFT_132__FPB_n345(net479_c1,net479);
INTERCONNECT SplitCLK_4_131_SplitCLK_0_129(net480_c1,net480);
INTERCONNECT SplitCLK_4_131_SplitCLK_4_130(net481_c1,net481);
INTERCONNECT SplitCLK_4_130_NOTT_64_n94(net482_c1,net482);
INTERCONNECT SplitCLK_4_130_DFFT_72__FBL_n285(net483_c1,net483);
INTERCONNECT SplitCLK_0_129_DFFT_133__FPB_n346(net484_c1,net484);
INTERCONNECT SplitCLK_0_129_DFFT_134__FPB_n347(net485_c1,net485);
INTERCONNECT GCLK_Pad_SplitCLK_0_255(GCLK_Pad,net486);

endmodule
