module TAP_route(
input GCLK_Pad,
input TMS_Pad,
output TDO_Pad,
output St_obs0_Pad,
output St_obs1_Pad,
output St_obs2_Pad);

wire net0_c1;
wire TDO_Pad;
wire TMS_Pad;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire St_obs0_Pad;
wire net275_c1;
wire St_obs1_Pad;
wire net276_c1;
wire St_obs2_Pad;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire net486_c1;
wire net486;
wire net487_c1;
wire net487;
wire net488_c1;
wire net488;
wire net489_c1;
wire net489;
wire net490_c1;
wire net490;
wire net491_c1;
wire net491;
wire net492_c1;
wire net492;
wire net493_c1;
wire net493;
wire net494_c1;
wire net494;
wire net495_c1;
wire net495;
wire net496_c1;
wire net496;
wire net497_c1;
wire net497;
wire net498_c1;
wire net498;
wire net499_c1;
wire net499;
wire net500_c1;
wire net500;
wire net501_c1;
wire net501;
wire net502_c1;
wire net502;
wire net503_c1;
wire net503;
wire net504_c1;
wire net504;
wire net505_c1;
wire net505;
wire net506_c1;
wire net506;
wire net507_c1;
wire net507;
wire net508_c1;
wire net508;
wire net509_c1;
wire net509;
wire net510_c1;
wire net510;
wire net511_c1;
wire net511;
wire net512_c1;
wire net512;
wire net513_c1;
wire net513;
wire net514_c1;
wire net514;
wire net515_c1;
wire net515;
wire net516_c1;
wire net516;
wire net517_c1;
wire net517;
wire net518_c1;
wire net518;
wire net519_c1;
wire net519;
wire net520_c1;
wire net520;
wire net521_c1;
wire net521;
wire net522_c1;
wire net522;
wire net523_c1;
wire net523;
wire net524_c1;
wire net524;
wire net525_c1;
wire net525;
wire net526_c1;
wire net526;
wire net527_c1;
wire net527;
wire net528_c1;
wire net528;
wire net529_c1;
wire net529;
wire net530_c1;
wire net530;
wire net531_c1;
wire net531;
wire net532_c1;
wire net532;
wire net533_c1;
wire net533;
wire net534_c1;
wire net534;
wire net535_c1;
wire net535;
wire net536_c1;
wire net536;
wire net537_c1;
wire net537;
wire net538_c1;
wire net538;
wire net539_c1;
wire net539;
wire net540_c1;
wire net540;
wire net541_c1;
wire net541;
wire net542_c1;
wire net542;
wire net543_c1;
wire net543;
wire net544_c1;
wire net544;
wire net545_c1;
wire net545;
wire net546_c1;
wire net546;
wire net547_c1;
wire net547;
wire net548_c1;
wire net548;
wire net549_c1;
wire net549;
wire net550_c1;
wire net550;
wire net551_c1;
wire net551;
wire net552_c1;
wire net552;
wire net553_c1;
wire net553;
wire net554_c1;
wire net554;
wire net555_c1;
wire net555;
wire net556_c1;
wire net556;
wire net557_c1;
wire net557;
wire net558_c1;
wire net558;
wire net559_c1;
wire net559;
wire net560_c1;
wire net560;
wire net561_c1;
wire net561;
wire net562_c1;
wire net562;
wire net563_c1;
wire net563;
wire net564_c1;
wire net564;
wire net565_c1;
wire net565;
wire net566_c1;
wire net566;
wire net567_c1;
wire net567;
wire net568_c1;
wire net568;
wire net569_c1;
wire net569;
wire net570_c1;
wire net570;
wire net571_c1;
wire net571;
wire net572_c1;
wire net572;
wire net573_c1;
wire net573;
wire net574_c1;
wire net574;
wire net575_c1;
wire net575;
wire net576_c1;
wire net576;
wire net577_c1;
wire net577;
wire net578_c1;
wire net578;
wire net579_c1;
wire net579;
wire net580_c1;
wire net580;
wire net581_c1;
wire net581;
wire net582_c1;
wire net582;
wire net583_c1;
wire net583;
wire net584_c1;
wire net584;
wire net585_c1;
wire net585;
wire net586_c1;
wire net586;
wire net587_c1;
wire net587;
wire net588_c1;
wire net588;
wire net589_c1;
wire net589;
wire net590_c1;
wire net590;
wire net591_c1;
wire net591;
wire net592_c1;
wire net592;
wire net593_c1;
wire net593;
wire net594_c1;
wire net594;
wire net595_c1;
wire net595;
wire net596_c1;
wire net596;
wire net597_c1;
wire net597;
wire net598_c1;
wire net598;
wire net599_c1;
wire net599;
wire net600_c1;
wire net600;
wire net601_c1;
wire net601;
wire net602_c1;
wire net602;
wire net603_c1;
wire net603;
wire net604_c1;
wire net604;
wire net605_c1;
wire net605;
wire net606_c1;
wire net606;
wire net607_c1;
wire net607;
wire net608_c1;
wire net608;
wire net609_c1;
wire net609;
wire net610_c1;
wire net610;
wire net611_c1;
wire net611;
wire net612_c1;
wire net612;
wire net613_c1;
wire net613;
wire net614_c1;
wire net614;
wire net615_c1;
wire net615;
wire net616_c1;
wire net616;
wire net617_c1;
wire net617;
wire net618_c1;
wire net618;
wire net619_c1;
wire net619;
wire net620_c1;
wire net620;
wire net621_c1;
wire net621;
wire net622_c1;
wire net622;
wire net623_c1;
wire net623;
wire net624_c1;
wire net624;
wire net625_c1;
wire net625;
wire net626_c1;
wire net626;
wire net627_c1;
wire net627;
wire net628_c1;
wire net628;
wire net629_c1;
wire net629;
wire net630_c1;
wire net630;
wire net631_c1;
wire net631;
wire net632_c1;
wire net632;
wire net633_c1;
wire net633;
wire net634_c1;
wire net634;
wire net635_c1;
wire net635;
wire net636_c1;
wire net636;
wire net637_c1;
wire net637;
wire net638_c1;
wire net638;
wire net639_c1;
wire net639;
wire net640_c1;
wire net640;
wire net641_c1;
wire net641;
wire net642_c1;
wire net642;
wire net643_c1;
wire net643;
wire net644_c1;
wire net644;
wire net645_c1;
wire net645;
wire net646_c1;
wire net646;
wire net647_c1;
wire net647;
wire net648_c1;
wire net648;
wire net649_c1;
wire net649;
wire net650_c1;
wire net650;
wire net651_c1;
wire net651;
wire net652_c1;
wire net652;
wire net653_c1;
wire net653;
wire net654_c1;
wire net654;
wire net655_c1;
wire net655;
wire net656_c1;
wire net656;
wire net657_c1;
wire net657;
wire net658_c1;
wire net658;
wire net659_c1;
wire net659;
wire net660_c1;
wire net660;
wire net661_c1;
wire net661;
wire net662_c1;
wire net662;
wire net663_c1;
wire net663;
wire net664_c1;
wire net664;
wire net665_c1;
wire net665;
wire net666_c1;
wire net666;
wire net667_c1;
wire net667;
wire net668_c1;
wire net668;
wire net669_c1;
wire net669;
wire net670_c1;
wire net670;
wire net671_c1;
wire net671;
wire net672_c1;
wire net672;
wire net673_c1;
wire net673;
wire net674_c1;
wire net674;
wire net675_c1;
wire net675;
wire net676_c1;
wire net676;
wire net677_c1;
wire net677;
wire net678_c1;
wire net678;
wire net679_c1;
wire net679;
wire net680_c1;
wire net680;
wire net681_c1;
wire net681;
wire net682_c1;
wire net682;
wire net683_c1;
wire net683;
wire net684_c1;
wire net684;
wire net685_c1;
wire net685;
wire net686_c1;
wire net686;
wire net687_c1;
wire net687;
wire net688_c1;
wire net688;
wire net689_c1;
wire net689;
wire net690_c1;
wire net690;
wire net691_c1;
wire net691;
wire net692_c1;
wire net692;
wire net693_c1;
wire net693;
wire net694_c1;
wire net694;
wire net695_c1;
wire net695;
wire net696_c1;
wire net696;
wire net697_c1;
wire net697;
wire net698_c1;
wire net698;
wire net699_c1;
wire net699;
wire net700_c1;
wire net700;
wire net701_c1;
wire net701;
wire net702_c1;
wire net702;
wire net703_c1;
wire net703;
wire net704_c1;
wire net704;
wire net705_c1;
wire net705;
wire net706_c1;
wire net706;
wire net707_c1;
wire net707;
wire net708_c1;
wire net708;
wire net709_c1;
wire net709;
wire net710_c1;
wire net710;
wire net711_c1;
wire net711;
wire net712_c1;
wire net712;
wire net713_c1;
wire net713;
wire net714_c1;
wire net714;
wire net715_c1;
wire net715;
wire net716_c1;
wire net716;
wire net717_c1;
wire net717;
wire net718_c1;
wire net718;
wire net719_c1;
wire net719;
wire net720_c1;
wire net720;
wire net721_c1;
wire net721;
wire net722_c1;
wire net722;
wire net723_c1;
wire net723;
wire net724_c1;
wire net724;
wire net725_c1;
wire net725;
wire net726_c1;
wire net726;
wire net727_c1;
wire net727;
wire net728_c1;
wire net728;
wire net729_c1;
wire net729;
wire net730_c1;
wire net730;
wire net731_c1;
wire net731;
wire net732_c1;
wire net732;
wire net733_c1;
wire net733;
wire net734_c1;
wire net734;
wire net735_c1;
wire net735;
wire net736_c1;
wire net736;
wire net737_c1;
wire net737;
wire net738_c1;
wire net738;
wire net739_c1;
wire net739;
wire net740_c1;
wire net740;
wire net741_c1;
wire net741;
wire net742_c1;
wire net742;
wire net743_c1;
wire net743;
wire net744_c1;
wire net744;
wire net745_c1;
wire net745;
wire net746_c1;
wire net746;
wire net747_c1;
wire net747;
wire net748_c1;
wire net748;
wire net749_c1;
wire net749;
wire net750_c1;
wire net750;
wire net751_c1;
wire net751;
wire net752_c1;
wire net752;
wire net753_c1;
wire net753;
wire net754_c1;
wire net754;
wire net755_c1;
wire net755;
wire net756_c1;
wire net756;
wire net757_c1;
wire net757;
wire net758_c1;
wire net758;
wire net759_c1;
wire net759;
wire net760_c1;
wire net760;
wire net761_c1;
wire net761;
wire net762_c1;
wire net762;
wire net763_c1;
wire net763;
wire net764_c1;
wire net764;
wire net765_c1;
wire net765;
wire net766_c1;
wire net766;
wire net767_c1;
wire net767;
wire net768_c1;
wire net768;
wire net769_c1;
wire net769;
wire net770_c1;
wire net770;
wire net771_c1;
wire net771;
wire net772_c1;
wire net772;
wire net773_c1;
wire net773;
wire net774_c1;
wire net774;
wire net775_c1;
wire net775;
wire net776_c1;
wire net776;
wire net777_c1;
wire net777;
wire net778_c1;
wire net778;
wire net779_c1;
wire net779;
wire net780_c1;
wire net780;
wire net781_c1;
wire net781;
wire net782_c1;
wire net782;
wire net783_c1;
wire net783;
wire net784_c1;
wire net784;
wire net785_c1;
wire net785;
wire net786_c1;
wire net786;
wire net787_c1;
wire net787;
wire net788_c1;
wire net788;
wire net789_c1;
wire net789;
wire net790_c1;
wire net790;
wire net791_c1;
wire net791;
wire net792_c1;
wire net792;
wire net793_c1;
wire net793;
wire net794_c1;
wire net794;
wire net795_c1;
wire net795;
wire net796_c1;
wire net796;
wire net797_c1;
wire net797;
wire net798_c1;
wire net798;
wire net799_c1;
wire net799;
wire net800_c1;
wire net800;
wire net801_c1;
wire net801;
wire net802_c1;
wire net802;
wire net803_c1;
wire net803;
wire net804_c1;
wire net804;
wire net805_c1;
wire net805;
wire net806_c1;
wire net806;
wire net807_c1;
wire net807;
wire net808_c1;
wire net808;
wire net809_c1;
wire net809;
wire net810_c1;
wire net810;
wire net811_c1;
wire net811;
wire net812_c1;
wire net812;
wire GCLK_Pad;
wire net813;
wire net814_c1;
wire net814;

XOR2T XOR2T_20_n32(net507,net153,net299,net9_c1);
AND2T AND2T_9_n21(net436,net248,net224,net3_c1);
DFFT DFFT_190_St_obs1(net493,net342,net275_c1);
NOTT NOTT_7_n19(net469,net245,net22_c1);
NOTT NOTT_8_n20(net470,net226,net2_c1);
DFFT DFFT_184_St_obs0(net435,net351,net274_c1);
DFFT DFFT_196_St_obs2(net645,net364,net276_c1);
AND2T AND2T_12_n24(net497,net268,net238,net10_c1);
AND2T AND2T_21_n33(net434,net157,net173,net12_c1);
AND2T AND2T_13_n25(net433,net218,net201,net13_c1);
AND2T AND2T_30_n42(net479,net158,net292,net15_c1);
AND2T AND2T_22_n34(net432,net115,net303,net16_c1);
AND2T AND2T_14_n26(net431,net180,net287,net17_c1);
AND2T AND2T_31_n43(net551,net211,net295,net19_c1);
AND2T AND2T_23_n35(net667,net244,net307,net20_c1);
AND2T AND2T_15_n27(net515,net141,net159,net21_c1);
AND2T AND2T_40_n52(net541,net223,net322,net24_c1);
AND2T AND2T_16_n28(net671,net258,net289,net27_c1);
AND2T AND2T_41_n53(net519,net262,net209,net29_c1);
AND2T AND2T_33_n45(net609,net25,net306,net30_c1);
AND2T AND2T_25_n37(net661,net205,net312,net31_c1);
AND2T AND2T_17_n29(net430,net272,net293,net32_c1);
AND2T AND2T_18_n30(net668,net135,net296,net4_c1);
AND2T AND2T_34_n46(net429,net97,net169,net36_c1);
AND2T AND2T_26_n38(net428,net31,net195,net37_c1);
AND2T AND2T_19_n31(net427,net186,net9,net6_c1);
AND2T AND2T_43_n55(net426,net203,net298,net40_c1);
AND2T AND2T_35_n47(net552,net125,net130,net41_c1);
AND2T AND2T_44_n56(net672,net156,net302,net46_c1);
AND2T AND2T_61_n73(net597,net188,net134,net49_c1);
AND2T AND2T_45_n57(net529,net207,net119,net51_c1);
AND2T AND2T_38_n50(net555,net52,net47,net14_c1);
AND2T AND2T_70_n82(net775,net213,net107,net54_c1);
AND2T AND2T_62_n74(net779,net194,net326,net55_c1);
AND2T AND2T_54_n66(net425,net50,net304,net56_c1);
AND2T AND2T_46_n58(net424,net234,net269,net57_c1);
AND2T AND2T_63_n75(net780,net99,net198,net60_c1);
AND2T AND2T_55_n67(net516,net229,net66,net61_c1);
AND2T AND2T_48_n60(net751,net212,net321,net23_c1);
AND2T AND2T_64_n76(net423,net60,net331,net65_c1);
AND2T AND2T_56_n68(net422,net265,net282,net66_c1);
AND2T AND2T_81_n93(net703,net192,net340,net67_c1);
AND2T AND2T_58_n70(net587,net187,net172,net33_c1);
AND2T AND2T_74_n86(net421,net98,net75,net72_c1);
AND2T AND2T_59_n71(net591,net221,net320,net38_c1);
AND2T AND2T_75_n87(net739,net147,net139,net75_c1);
AND2T AND2T_84_n96(net752,net271,net345,net77_c1);
AND2T AND2T_69_n81(net785,net230,net310,net48_c1);
AND2T AND2T_85_n97(net420,net133,net353,net79_c1);
AND2T AND2T_79_n91(net461,net63,net330,net58_c1);
AND2T AND2T_87_n99(net789,net106,net329,net82_c1);
OR2T OR2T_32_n44(net563,net189,net247,net25_c1);
OR2T OR2T_50_n62(net619,net28,net18,net34_c1);
OR2T OR2T_42_n54(net419,net29,net24,net35_c1);
OR2T OR2T_51_n63(net418,net34,net327,net39_c1);
OR2T OR2T_27_n39(net483,net202,net190,net42_c1);
OR2T OR2T_28_n40(net588,net42,net317,net8_c1);
OR2T OR2T_60_n72(net601,net191,net273,net44_c1);
OR2T OR2T_52_n64(net417,net100,net101,net45_c1);
OR2T OR2T_36_n48(net610,net199,net193,net47_c1);
OR2T OR2T_29_n41(net416,net8,net291,net11_c1);
OR2T OR2T_53_n65(net761,net216,net124,net50_c1);
OR2T OR2T_37_n49(net545,net111,net316,net52_c1);
OR2T OR2T_39_n51(net415,net14,net30,net18_c1);
OR2T OR2T_71_n83(net733,net104,net183,net59_c1);
OR2T OR2T_47_n59(net662,net51,net305,net62_c1);
OR2T OR2T_80_n92(net414,net252,net140,net63_c1);
OR2T OR2T_72_n84(net413,net59,net315,net64_c1);
OR2T OR2T_49_n61(net412,net23,net40,net28_c1);
OR2T OR2T_73_n85(net556,net129,net113,net68_c1);
OR2T OR2T_65_n77(net786,net200,net55,net69_c1);
OR2T OR2T_57_n69(net484,net114,net311,net70_c1);
OR2T OR2T_82_n94(net704,net67,net58,net71_c1);
OR2T OR2T_66_n78(net411,net69,net44,net73_c1);
DFFT DFFT_178_TDO(net410,net359,net0_c1);
OR2T OR2T_83_n95(net707,net71,net109,net74_c1);
OR2T OR2T_67_n79(net409,net73,net341,net76_c1);
OR2T OR2T_68_n80(net530,net76,net346,net43_c1);
OR2T OR2T_76_n88(net734,net103,net319,net78_c1);
OR2T OR2T_77_n89(net602,net78,net68,net80_c1);
OR2T OR2T_78_n90(net729,net80,net325,net53_c1);
OR2T OR2T_86_n98(net743,net79,net77,net81_c1);
NOTT NOTT_10_n22(net451,net260,net5_c1);
NOTT NOTT_11_n23(net452,net246,net7_c1);
NOTT NOTT_24_n36(net408,net254,net26_c1);
AND2T AND2T_92_n104(net407,net241,net261,net87_c1);
AND2T AND2T_93_n105(net503,net152,net171,net89_c1);
AND2T AND2T_94_n106(net504,net270,net257,net91_c1);
AND2T AND2T_95_n113(net406,net164,net22,net88_c1);
AND2T AND2T_88_n100(net797,net196,net336,net83_c1);
AND2T AND2T_96_n114(net405,net266,net5,net90_c1);
AND2T AND2T_97_n115(net649,net277,net283,net93_c1);
DFFT DFFT_101__FPB_n128(net623,net138,net286_c1);
DFFT DFFT_110__FBL_n392(net404,net367,net279_c1);
DFFT DFFT_102__FPB_n129(net755,net231,net288_c1);
DFFT DFFT_111__FBL_n393(net403,net368,net280_c1);
DFFT DFFT_103__FBL_n385(net473,net39,net281_c1);
DFFT DFFT_104__FBL_n386(net525,net204,net282_c1);
DFFT DFFT_120__FPB_n402(net402,net168,net290_c1);
DFFT DFFT_112__FPB_n394(net401,net222,net356_c1);
DFFT DFFT_105__FBL_n387(net400,net356,net283_c1);
DFFT DFFT_121__FPB_n403(net801,net290,net293_c1);
DFFT DFFT_113__FPB_n395(net695,net233,net360_c1);
DFFT DFFT_106__FBL_n388(net696,net360,net284_c1);
DFFT DFFT_130__FPB_n412(net546,net151,net295_c1);
DFFT DFFT_122__FPB_n404(net657,net232,net296_c1);
DFFT DFFT_114__FPB_n396(net685,net145,net363_c1);
DFFT DFFT_107__FBL_n389(net399,net112,net285_c1);
DFFT DFFT_131__FPB_n413(net613,net120,net297_c1);
DFFT DFFT_123__FPB_n405(net508,net251,net299_c1);
DFFT DFFT_115__FPB_n397(net398,net227,net366_c1);
DFFT DFFT_108__FBL_n390(net397,net363,net277_c1);
DFFT DFFT_140__FPB_n422(net717,net259,net302_c1);
DFFT DFFT_132__FPB_n414(net614,net297,net301_c1);
DFFT DFFT_124__FPB_n406(net542,net237,net303_c1);
DFFT DFFT_116__FPB_n398(net686,net132,net367_c1);
DFFT DFFT_109__FBL_n391(net639,net366,net278_c1);
DFFT DFFT_141__FPB_n423(net730,net57,net305_c1);
DFFT DFFT_133__FPB_n415(net396,net301,net306_c1);
DFFT DFFT_125__FPB_n407(net395,net144,net307_c1);
DFFT DFFT_117__FPB_n399(net640,net217,net368_c1);
DFFT DFFT_118__FPB_n400(net498,net178,net287_c1);
DFFT DFFT_150__FPB_n432(net526,net61,net311_c1);
DFFT DFFT_142__FPB_n424(net394,net210,net308_c1);
DFFT DFFT_134__FPB_n416(net564,net215,net309_c1);
DFFT DFFT_126__FPB_n408(net658,net162,net312_c1);
DFFT DFFT_119__FPB_n401(net740,net179,net289_c1);
DFFT DFFT_151__FPB_n433(net765,net122,net313_c1);
DFFT DFFT_143__FPB_n425(net393,net308,net314_c1);
DFFT DFFT_135__FPB_n417(net392,net309,net316_c1);
DFFT DFFT_127__FPB_n409(net391,net6,net317_c1);
OR2T OR2T_90_n102(net798,net84,net81,net85_c1);
OR2T OR2T_91_n103(net713,net85,net339,net86_c1);
DFFT DFFT_128__FPB_n410(net390,net184,net291_c1);
DFFT DFFT_160__FPB_n442(net598,net72,net319_c1);
DFFT DFFT_152__FPB_n434(net762,net313,net320_c1);
DFFT DFFT_144__FPB_n426(net624,net314,net321_c1);
DFFT DFFT_136__FPB_n418(net389,net267,net322_c1);
OR2T OR2T_89_n101(net807,net83,net82,net84_c1);
DFFT DFFT_129__FPB_n411(net474,net163,net292_c1);
DFFT DFFT_161__FPB_n443(net388,net64,net325_c1);
DFFT DFFT_153__FPB_n435(net387,net110,net326_c1);
DFFT DFFT_145__FPB_n427(net592,net11,net327_c1);
DFFT DFFT_137__FPB_n419(net386,net127,net324_c1);
DFFT DFFT_138__FPB_n420(net573,net324,net294_c1);
DFFT DFFT_170__FPB_n452(net766,net323,net329_c1);
DFFT DFFT_162__FPB_n444(net462,net12,net330_c1);
DFFT DFFT_154__FPB_n436(net385,net118,net331_c1);
DFFT DFFT_146__FPB_n428(net802,net236,net328_c1);
DFFT DFFT_139__FPB_n421(net574,net294,net298_c1);
DFFT DFFT_171__FPB_n453(net790,net208,net336_c1);
DFFT DFFT_163__FPB_n445(net714,net255,net333_c1);
DFFT DFFT_155__FPB_n437(net384,net70,net334_c1);
DFFT DFFT_147__FPB_n429(net383,net328,net335_c1);
DFFT DFFT_148__FPB_n430(net811,net335,net300_c1);
DFFT DFFT_180__FPB_n462(net457,net332,net338_c1);
DFFT DFFT_172__FPB_n454(net708,net74,net339_c1);
DFFT DFFT_164__FPB_n446(net382,net333,net340_c1);
DFFT DFFT_156__FPB_n438(net520,net334,net341_c1);
DFFT DFFT_149__FPB_n431(net812,net300,net304_c1);
DFFT DFFT_181__FPB_n463(net458,net338,net343_c1);
DFFT DFFT_173__FPB_n455(net381,net155,net344_c1);
DFFT DFFT_165__FPB_n447(net744,net123,net345_c1);
DFFT DFFT_157__FPB_n439(net620,net56,net346_c1);
DFFT DFFT_158__FPB_n440(net718,net170,net310_c1);
DFFT DFFT_182__FPB_n464(net380,net343,net347_c1);
DFFT DFFT_174__FPB_n456(net577,net344,net348_c1);
DFFT DFFT_166__FPB_n448(net379,net143,net349_c1);
SPLITT Split_200_n482(net2,net150_c1,net242_c1);
SPLITT Split_201_n483(net242,net158_c1,net248_c1);
SPLITT Split_202_n484(net150,net164_c1,net252_c1);
SPLITT Split_210_n492(net17,net161_c1,net253_c1);
SPLITT Split_203_n485(net3,net167_c1,net257_c1);
SPLITT Split_211_n493(net253,net169_c1,net258_c1);
SPLITT Split_220_n502(net96,net98_c1,net188_c1);
SPLITT Split_204_n486(net167,net171_c1,net261_c1);
SPLITT Split_212_n494(net161,net172_c1,net262_c1);
SPLITT Split_221_n503(net16,net101_c1,net190_c1);
SPLITT Split_205_n487(net7,net177_c1,net266_c1);
SPLITT Split_213_n495(net21,net176_c1,net267_c1);
SPLITT Split_222_n504(net20,net102_c1,net192_c1);
SPLITT Split_230_n512(net36,net104_c1,net193_c1);
SPLITT Split_206_n488(net177,net180_c1,net268_c1);
SPLITT Split_214_n496(net176,net179_c1,net269_c1);
SPLITT Split_223_n505(net102,net107_c1,net195_c1);
SPLITT Split_231_n513(net41,net105_c1,net196_c1);
SPLITT Split_207_n489(net10,net181_c1,net270_c1);
SPLITT Split_215_n497(net27,net182_c1,net271_c1);
SPLITT Split_224_n506(net26,net110_c1,net198_c1);
SPLITT Split_232_n514(net105,net111_c1,net199_c1);
SPLITT Split_240_n522(net65,net109_c1,net200_c1);
SPLITT Split_208_n490(net181,net152_c1,net241_c1);
SPLITT Split_216_n498(net182,net183_c1,net272_c1);
SPLITT Split_225_n507(net37,net114_c1,net202_c1);
SPLITT Split_233_n515(net35,net113_c1,net203_c1);
SPLITT Split_241_n523(net43,net112_c1,net204_c1);
SPLITT Split_209_n491(net13,net155_c1,net247_c1);
SPLITT Split_217_n499(net32,net184_c1,net273_c1);
SPLITT Split_218_n500(net4,net96_c1,net185_c1);
SPLITT Split_226_n508(net15,net116_c1,net206_c1);
SPLITT Split_234_n516(net46,net118_c1,net207_c1);
SPLITT Split_242_n524(net48,net117_c1,net208_c1);
SPLITT Split_250_n532(net108,net119_c1,net209_c1);
SPLITT Split_219_n501(net185,net97_c1,net186_c1);
SPLITT Split_227_n509(net206,net125_c1,net211_c1);
SPLITT Split_235_n517(net62,net124_c1,net212_c1);
SPLITT Split_243_n525(net117,net123_c1,net213_c1);
SPLITT Split_251_n533(net90,net121_c1,net214_c1);
SPLITT Split_228_n510(net116,net99_c1,net187_c1);
SPLITT Split_236_n518(net45,net129_c1,net216_c1);
SPLITT Split_244_n526(net53,net128_c1,net217_c1);
SPLITT Split_252_n534(net214,net130_c1,net218_c1);
SPLITT Split_260_n542(net92,net126_c1,net219_c1);
SPLITT Split_229_n511(net19,net100_c1,net189_c1);
SPLITT Split_237_n519(net33,net133_c1,net221_c1);
SPLITT Split_245_n527(net128,net132_c1,net222_c1);
SPLITT Split_253_n535(net121,net134_c1,net223_c1);
SPLITT Split_261_n543(net219,net135_c1,net224_c1);
SPLITT Split_238_n520(net38,net103_c1,net191_c1);
SPLITT Split_246_n528(net86,net137_c1,net227_c1);
SPLITT Split_254_n536(net93,net136_c1,net228_c1);
SPLITT Split_262_n544(net126,net140_c1,net229_c1);
SPLITT Split_270_n552(net220,net139_c1,net230_c1);
SPLITT Split_239_n521(net49,net106_c1,net194_c1);
SPLITT Split_247_n529(net137,net145_c1,net233_c1);
SPLITT Split_255_n537(net228,net147_c1,net234_c1);
SPLITT Split_263_n545(net94,net142_c1,net235_c1);
SPLITT Split_271_n553(net131,net143_c1,net236_c1);
SPLITT Split_248_n530(net88,net108_c1,net197_c1);
SPLITT Split_256_n538(net136,net151_c1,net237_c1);
SPLITT Split_264_n546(net235,net153_c1,net238_c1);
SPLITT Split_272_n554(net281,net149_c1,net239_c1);
SPLITT Split_280_n562(net278,net148_c1,net240_c1);
SPLITT Split_249_n531(net197,net115_c1,net201_c1);
SPLITT Split_257_n539(net95,net154_c1,net243_c1);
SPLITT Split_265_n547(net142,net156_c1,net244_c1);
SPLITT Split_273_n555(net239,net159_c1,net245_c1);
SPLITT Split_281_n563(net240,net157_c1,net246_c1);
DFFT DFFT_159__FPB_n441(net776,net54,net315_c1);
SPLITT Split_258_n540(net243,net120_c1,net205_c1);
DFFT DFFT_191__FPB_n473(net691,net91,net350_c1);
DFFT DFFT_183__FPB_n465(net378,net347,net351_c1);
DFFT DFFT_175__FPB_n457(net578,net348,net352_c1);
DFFT DFFT_167__FPB_n449(net808,net349,net353_c1);
SPLITT Split_266_n548(net286,net160_c1,net249_c1);
SPLITT Split_274_n556(net149,net163_c1,net250_c1);
SPLITT Split_282_n564(net148,net162_c1,net251_c1);
SPLITT Split_259_n541(net154,net122_c1,net210_c1);
SPLITT Split_267_n549(net249,net168_c1,net254_c1);
SPLITT Split_275_n557(net284,net166_c1,net255_c1);
SPLITT Split_283_n565(net280,net165_c1,net256_c1);
SPLITT Split_268_n550(net160,net127_c1,net215_c1);
SPLITT Split_276_n558(net166,net170_c1,net259_c1);
SPLITT Split_284_n566(net256,net173_c1,net260_c1);
SPLITT Split_269_n551(net288,net131_c1,net220_c1);
SPLITT Split_197_n479(net1,net175_c1,net263_c1);
SPLITT Split_277_n559(net285,net174_c1,net264_c1);
SPLITT Split_285_n567(net165,net178_c1,net265_c1);
SPLITT Split_198_n480(net263,net138_c1,net225_c1);
SPLITT Split_278_n560(net264,net141_c1,net226_c1);
SPLITT Split_199_n481(net175,net146_c1,net231_c1);
SPLITT Split_279_n561(net174,net144_c1,net232_c1);
NOTT NOTT_100_n124(net650,net814,net94_c1);
DFFT DFFT_168__FPB_n450(net756,net146,net318_c1);
DFFT DFFT_192__FPB_n474(net692,net350,net354_c1);
DFFT DFFT_176__FPB_n458(net567,net352,net355_c1);
DFFT DFFT_169__FPB_n451(net377,net318,net323_c1);
DFFT DFFT_193__FPB_n475(net681,net354,net357_c1);
DFFT DFFT_185__FPB_n467(net376,net89,net358_c1);
DFFT DFFT_177__FPB_n459(net568,net355,net359_c1);
DFFT DFFT_194__FPB_n476(net682,net357,net361_c1);
DFFT DFFT_186__FPB_n468(net375,net358,net362_c1);
DFFT DFFT_179__FPB_n461(net374,net87,net332_c1);
DFFT DFFT_195__FPB_n477(net373,net361,net364_c1);
DFFT DFFT_187__FPB_n469(net372,net362,net365_c1);
DFFT DFFT_188__FPB_n470(net646,net365,net337_c1);
NOTT NOTT_98_n116(net371,net225,net95_c1);
NOTT NOTT_99_n123(net480,net250,net92_c1);
DFFT DFFT_189__FPB_n471(net494,net337,net342_c1);
SPLITT SplitCLK_4_191(net810,net811_c1,net812_c1);
SPLITT SplitCLK_0_192(net803,net809_c1,net810_c1);
SPLITT SplitCLK_4_193(net806,net807_c1,net808_c1);
SPLITT SplitCLK_2_194(net804,net805_c1,net806_c1);
SPLITT SplitCLK_4_195(net791,net804_c1,net803_c1);
SPLITT SplitCLK_4_196(net800,net802_c1,net801_c1);
SPLITT SplitCLK_6_197(net793,net800_c1,net799_c1);
SPLITT SplitCLK_4_198(net796,net798_c1,net797_c1);
SPLITT SplitCLK_2_199(net794,net796_c1,net795_c1);
SPLITT SplitCLK_6_200(net792,net793_c1,net794_c1);
SPLITT SplitCLK_6_201(net767,net791_c1,net792_c1);
SPLITT SplitCLK_4_202(net788,net789_c1,net790_c1);
SPLITT SplitCLK_6_203(net781,net788_c1,net787_c1);
SPLITT SplitCLK_4_204(net784,net786_c1,net785_c1);
SPLITT SplitCLK_4_205(net782,net783_c1,net784_c1);
SPLITT SplitCLK_0_206(net769,net781_c1,net782_c1);
SPLITT SplitCLK_4_207(net778,net780_c1,net779_c1);
SPLITT SplitCLK_6_208(net771,net778_c1,net777_c1);
SPLITT SplitCLK_4_209(net774,net776_c1,net775_c1);
SPLITT SplitCLK_6_210(net772,net774_c1,net773_c1);
SPLITT SplitCLK_4_211(net770,net772_c1,net771_c1);
SPLITT SplitCLK_4_212(net768,net770_c1,net769_c1);
SPLITT SplitCLK_0_213(net719,net767_c1,net768_c1);
SPLITT SplitCLK_4_214(net764,net765_c1,net766_c1);
SPLITT SplitCLK_2_215(net757,net763_c1,net764_c1);
SPLITT SplitCLK_4_216(net760,net761_c1,net762_c1);
SPLITT SplitCLK_4_217(net758,net759_c1,net760_c1);
SPLITT SplitCLK_0_218(net745,net757_c1,net758_c1);
SPLITT SplitCLK_0_219(net754,net755_c1,net756_c1);
SPLITT SplitCLK_2_220(net747,net753_c1,net754_c1);
SPLITT SplitCLK_4_221(net750,net752_c1,net751_c1);
SPLITT SplitCLK_4_222(net748,net749_c1,net750_c1);
SPLITT SplitCLK_2_223(net746,net748_c1,net747_c1);
SPLITT SplitCLK_6_224(net721,net745_c1,net746_c1);
SPLITT SplitCLK_4_225(net742,net743_c1,net744_c1);
SPLITT SplitCLK_2_226(net735,net741_c1,net742_c1);
SPLITT SplitCLK_4_227(net738,net740_c1,net739_c1);
SPLITT SplitCLK_2_228(net736,net737_c1,net738_c1);
SPLITT SplitCLK_4_229(net723,net736_c1,net735_c1);
SPLITT SplitCLK_4_230(net732,net734_c1,net733_c1);
SPLITT SplitCLK_2_231(net725,net732_c1,net731_c1);
SPLITT SplitCLK_4_232(net728,net730_c1,net729_c1);
SPLITT SplitCLK_4_233(net726,net727_c1,net728_c1);
SPLITT SplitCLK_2_234(net724,net726_c1,net725_c1);
SPLITT SplitCLK_4_235(net722,net724_c1,net723_c1);
SPLITT SplitCLK_2_236(net720,net722_c1,net721_c1);
SPLITT SplitCLK_6_237(net625,net719_c1,net720_c1);
SPLITT SplitCLK_4_238(net716,net717_c1,net718_c1);
SPLITT SplitCLK_6_239(net709,net716_c1,net715_c1);
SPLITT SplitCLK_4_240(net712,net713_c1,net714_c1);
SPLITT SplitCLK_2_241(net710,net711_c1,net712_c1);
SPLITT SplitCLK_0_242(net697,net709_c1,net710_c1);
SPLITT SplitCLK_4_243(net706,net707_c1,net708_c1);
SPLITT SplitCLK_6_244(net699,net706_c1,net705_c1);
SPLITT SplitCLK_4_245(net702,net704_c1,net703_c1);
SPLITT SplitCLK_4_246(net700,net701_c1,net702_c1);
SPLITT SplitCLK_2_247(net698,net700_c1,net699_c1);
SPLITT SplitCLK_6_248(net673,net697_c1,net698_c1);
SPLITT SplitCLK_4_249(net694,net695_c1,net696_c1);
SPLITT SplitCLK_0_250(net687,net694_c1,net693_c1);
SPLITT SplitCLK_4_251(net690,net692_c1,net691_c1);
SPLITT SplitCLK_4_252(net688,net689_c1,net690_c1);
SPLITT SplitCLK_4_253(net675,net688_c1,net687_c1);
SPLITT SplitCLK_4_254(net684,net686_c1,net685_c1);
SPLITT SplitCLK_6_255(net677,net684_c1,net683_c1);
SPLITT SplitCLK_4_256(net680,net682_c1,net681_c1);
SPLITT SplitCLK_4_257(net678,net679_c1,net680_c1);
SPLITT SplitCLK_2_258(net676,net678_c1,net677_c1);
SPLITT SplitCLK_4_259(net674,net676_c1,net675_c1);
SPLITT SplitCLK_0_260(net627,net673_c1,net674_c1);
SPLITT SplitCLK_4_261(net670,net671_c1,net672_c1);
SPLITT SplitCLK_4_262(net663,net669_c1,net670_c1);
SPLITT SplitCLK_4_263(net666,net668_c1,net667_c1);
SPLITT SplitCLK_2_264(net664,net665_c1,net666_c1);
SPLITT SplitCLK_4_265(net651,net663_c1,net664_c1);
SPLITT SplitCLK_4_266(net660,net662_c1,net661_c1);
SPLITT SplitCLK_2_267(net653,net659_c1,net660_c1);
SPLITT SplitCLK_4_268(net656,net657_c1,net658_c1);
SPLITT SplitCLK_4_269(net654,net655_c1,net656_c1);
SPLITT SplitCLK_2_270(net652,net654_c1,net653_c1);
SPLITT SplitCLK_2_271(net629,net651_c1,net652_c1);
SPLITT SplitCLK_4_272(net648,net650_c1,net649_c1);
SPLITT SplitCLK_2_273(net641,net647_c1,net648_c1);
SPLITT SplitCLK_4_274(net644,net646_c1,net645_c1);
SPLITT SplitCLK_4_275(net642,net643_c1,net644_c1);
SPLITT SplitCLK_0_276(net631,net641_c1,net642_c1);
SPLITT SplitCLK_4_277(net638,net640_c1,net639_c1);
SPLITT SplitCLK_4_278(net633,net637_c1,net638_c1);
SPLITT SplitCLK_4_279(net634,net635_c1,net636_c1);
SPLITT SplitCLK_6_280(net632,net633_c1,net634_c1);
SPLITT SplitCLK_4_281(net630,net632_c1,net631_c1);
SPLITT SplitCLK_2_282(net628,net630_c1,net629_c1);
SPLITT SplitCLK_4_283(net626,net628_c1,net627_c1);
SPLITT SplitCLK_0_284(net369,net625_c1,net626_c1);
SPLITT SplitCLK_4_285(net622,net623_c1,net624_c1);
SPLITT SplitCLK_4_286(net615,net621_c1,net622_c1);
SPLITT SplitCLK_4_287(net618,net620_c1,net619_c1);
SPLITT SplitCLK_2_288(net616,net617_c1,net618_c1);
SPLITT SplitCLK_0_289(net603,net615_c1,net616_c1);
SPLITT SplitCLK_4_290(net612,net614_c1,net613_c1);
SPLITT SplitCLK_6_291(net605,net612_c1,net611_c1);
SPLITT SplitCLK_4_292(net608,net610_c1,net609_c1);
SPLITT SplitCLK_4_293(net606,net607_c1,net608_c1);
SPLITT SplitCLK_6_294(net604,net606_c1,net605_c1);
SPLITT SplitCLK_6_295(net579,net603_c1,net604_c1);
SPLITT SplitCLK_4_296(net600,net601_c1,net602_c1);
SPLITT SplitCLK_6_297(net593,net600_c1,net599_c1);
SPLITT SplitCLK_4_298(net596,net598_c1,net597_c1);
SPLITT SplitCLK_4_299(net594,net595_c1,net596_c1);
SPLITT SplitCLK_0_300(net581,net593_c1,net594_c1);
SPLITT SplitCLK_4_301(net590,net591_c1,net592_c1);
SPLITT SplitCLK_6_302(net583,net590_c1,net589_c1);
SPLITT SplitCLK_4_303(net586,net588_c1,net587_c1);
SPLITT SplitCLK_2_304(net584,net585_c1,net586_c1);
SPLITT SplitCLK_6_305(net582,net583_c1,net584_c1);
SPLITT SplitCLK_4_306(net580,net582_c1,net581_c1);
SPLITT SplitCLK_0_307(net531,net579_c1,net580_c1);
SPLITT SplitCLK_4_308(net576,net577_c1,net578_c1);
SPLITT SplitCLK_6_309(net569,net576_c1,net575_c1);
SPLITT SplitCLK_4_310(net572,net573_c1,net574_c1);
SPLITT SplitCLK_6_311(net570,net572_c1,net571_c1);
SPLITT SplitCLK_4_312(net557,net570_c1,net569_c1);
SPLITT SplitCLK_4_313(net566,net568_c1,net567_c1);
SPLITT SplitCLK_6_314(net559,net566_c1,net565_c1);
SPLITT SplitCLK_4_315(net562,net563_c1,net564_c1);
SPLITT SplitCLK_2_316(net560,net561_c1,net562_c1);
SPLITT SplitCLK_6_317(net558,net559_c1,net560_c1);
SPLITT SplitCLK_6_318(net533,net557_c1,net558_c1);
SPLITT SplitCLK_4_319(net554,net556_c1,net555_c1);
SPLITT SplitCLK_2_320(net547,net553_c1,net554_c1);
SPLITT SplitCLK_4_321(net550,net551_c1,net552_c1);
SPLITT SplitCLK_4_322(net548,net549_c1,net550_c1);
SPLITT SplitCLK_0_323(net535,net547_c1,net548_c1);
SPLITT SplitCLK_4_324(net544,net545_c1,net546_c1);
SPLITT SplitCLK_2_325(net537,net543_c1,net544_c1);
SPLITT SplitCLK_4_326(net540,net542_c1,net541_c1);
SPLITT SplitCLK_4_327(net538,net539_c1,net540_c1);
SPLITT SplitCLK_4_328(net536,net537_c1,net538_c1);
SPLITT SplitCLK_4_329(net534,net536_c1,net535_c1);
SPLITT SplitCLK_6_330(net532,net533_c1,net534_c1);
SPLITT SplitCLK_6_331(net437,net531_c1,net532_c1);
SPLITT SplitCLK_4_332(net528,net529_c1,net530_c1);
SPLITT SplitCLK_6_333(net521,net528_c1,net527_c1);
SPLITT SplitCLK_4_334(net524,net526_c1,net525_c1);
SPLITT SplitCLK_2_335(net522,net523_c1,net524_c1);
SPLITT SplitCLK_0_336(net509,net521_c1,net522_c1);
SPLITT SplitCLK_4_337(net518,net520_c1,net519_c1);
SPLITT SplitCLK_4_338(net511,net517_c1,net518_c1);
SPLITT SplitCLK_4_339(net514,net515_c1,net516_c1);
SPLITT SplitCLK_4_340(net512,net513_c1,net514_c1);
SPLITT SplitCLK_6_341(net510,net511_c1,net512_c1);
SPLITT SplitCLK_6_342(net485,net509_c1,net510_c1);
SPLITT SplitCLK_4_343(net506,net508_c1,net507_c1);
SPLITT SplitCLK_6_344(net499,net506_c1,net505_c1);
SPLITT SplitCLK_4_345(net502,net504_c1,net503_c1);
SPLITT SplitCLK_2_346(net500,net501_c1,net502_c1);
SPLITT SplitCLK_0_347(net487,net499_c1,net500_c1);
SPLITT SplitCLK_4_348(net496,net497_c1,net498_c1);
SPLITT SplitCLK_2_349(net489,net495_c1,net496_c1);
SPLITT SplitCLK_4_350(net492,net493_c1,net494_c1);
SPLITT SplitCLK_4_351(net490,net491_c1,net492_c1);
SPLITT SplitCLK_2_352(net488,net490_c1,net489_c1);
SPLITT SplitCLK_4_353(net486,net488_c1,net487_c1);
SPLITT SplitCLK_0_354(net439,net485_c1,net486_c1);
SPLITT SplitCLK_4_355(net482,net484_c1,net483_c1);
SPLITT SplitCLK_2_356(net475,net481_c1,net482_c1);
SPLITT SplitCLK_4_357(net478,net479_c1,net480_c1);
SPLITT SplitCLK_2_358(net476,net477_c1,net478_c1);
SPLITT SplitCLK_0_359(net463,net475_c1,net476_c1);
SPLITT SplitCLK_4_360(net472,net473_c1,net474_c1);
SPLITT SplitCLK_2_361(net465,net472_c1,net471_c1);
SPLITT SplitCLK_4_362(net468,net469_c1,net470_c1);
SPLITT SplitCLK_4_363(net466,net467_c1,net468_c1);
SPLITT SplitCLK_4_364(net464,net465_c1,net466_c1);
SPLITT SplitCLK_6_365(net441,net463_c1,net464_c1);
SPLITT SplitCLK_4_366(net460,net462_c1,net461_c1);
SPLITT SplitCLK_6_367(net453,net460_c1,net459_c1);
SPLITT SplitCLK_4_368(net456,net458_c1,net457_c1);
SPLITT SplitCLK_4_369(net454,net455_c1,net456_c1);
SPLITT SplitCLK_0_370(net443,net453_c1,net454_c1);
SPLITT SplitCLK_4_371(net450,net452_c1,net451_c1);
SPLITT SplitCLK_6_372(net445,net450_c1,net449_c1);
SPLITT SplitCLK_4_373(net446,net447_c1,net448_c1);
SPLITT SplitCLK_2_374(net444,net446_c1,net445_c1);
SPLITT SplitCLK_4_375(net442,net444_c1,net443_c1);
SPLITT SplitCLK_2_376(net440,net442_c1,net441_c1);
SPLITT SplitCLK_4_377(net438,net440_c1,net439_c1);
SPLITT SplitCLK_2_378(net370,net438_c1,net437_c1);
wire dummy0;
SPLITT SplitCLK_2_379(net523,net436_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_2_380(net447,net435_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_381(net459,net434_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_382(net539,net433_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_4_383(net549,net432_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_2_384(net495,net431_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_2_385(net731,net430_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_2_386(net705,net429_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_2_387(net669,net428_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_2_388(net659,net427_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_2_389(net553,net426_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_2_390(net795,net425_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_4_391(net773,net424_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_4_392(net783,net423_c1,dummy13);
wire dummy14;
SPLITT SplitCLK_2_393(net505,net422_c1,dummy14);
wire dummy15;
SPLITT SplitCLK_2_394(net727,net421_c1,dummy15);
wire dummy16;
SPLITT SplitCLK_4_395(net759,net420_c1,dummy16);
wire dummy17;
SPLITT SplitCLK_2_396(net481,net419_c1,dummy17);
wire dummy18;
SPLITT SplitCLK_2_397(net589,net418_c1,dummy18);
wire dummy19;
SPLITT SplitCLK_2_398(net543,net417_c1,dummy19);
wire dummy20;
SPLITT SplitCLK_2_399(net585,net416_c1,dummy20);
wire dummy21;
SPLITT SplitCLK_2_400(net617,net415_c1,dummy21);
wire dummy22;
SPLITT SplitCLK_2_401(net477,net414_c1,dummy22);
wire dummy23;
SPLITT SplitCLK_2_402(net741,net413_c1,dummy23);
wire dummy24;
SPLITT SplitCLK_2_403(net749,net412_c1,dummy24);
wire dummy25;
SPLITT SplitCLK_2_404(net595,net411_c1,dummy25);
wire dummy26;
SPLITT SplitCLK_2_405(net565,net410_c1,dummy26);
wire dummy27;
SPLITT SplitCLK_2_406(net527,net409_c1,dummy27);
wire dummy28;
SPLITT SplitCLK_2_407(net787,net408_c1,dummy28);
wire dummy29;
SPLITT SplitCLK_2_408(net501,net407_c1,dummy29);
wire dummy30;
SPLITT SplitCLK_2_409(net467,net406_c1,dummy30);
wire dummy31;
SPLITT SplitCLK_2_410(net449,net405_c1,dummy31);
wire dummy32;
SPLITT SplitCLK_2_411(net683,net404_c1,dummy32);
wire dummy33;
SPLITT SplitCLK_2_412(net637,net403_c1,dummy33);
wire dummy34;
SPLITT SplitCLK_2_413(net805,net402_c1,dummy34);
wire dummy35;
SPLITT SplitCLK_2_414(net689,net401_c1,dummy35);
wire dummy36;
SPLITT SplitCLK_4_415(net693,net400_c1,dummy36);
wire dummy37;
SPLITT SplitCLK_2_416(net655,net399_c1,dummy37);
wire dummy38;
SPLITT SplitCLK_2_417(net647,net398_c1,dummy38);
wire dummy39;
SPLITT SplitCLK_4_418(net701,net397_c1,dummy39);
wire dummy40;
SPLITT SplitCLK_2_419(net607,net396_c1,dummy40);
wire dummy41;
SPLITT SplitCLK_2_420(net665,net395_c1,dummy41);
wire dummy42;
SPLITT SplitCLK_2_421(net753,net394_c1,dummy42);
wire dummy43;
SPLITT SplitCLK_2_422(net621,net393_c1,dummy43);
wire dummy44;
SPLITT SplitCLK_2_423(net561,net392_c1,dummy44);
wire dummy45;
SPLITT SplitCLK_2_424(net513,net391_c1,dummy45);
wire dummy46;
SPLITT SplitCLK_2_425(net599,net390_c1,dummy46);
wire dummy47;
SPLITT SplitCLK_2_426(net471,net389_c1,dummy47);
wire dummy48;
SPLITT SplitCLK_2_427(net737,net388_c1,dummy48);
wire dummy49;
SPLITT SplitCLK_2_428(net777,net387_c1,dummy49);
wire dummy50;
SPLITT SplitCLK_2_429(net571,net386_c1,dummy50);
wire dummy51;
SPLITT SplitCLK_2_430(net715,net385_c1,dummy51);
wire dummy52;
SPLITT SplitCLK_2_431(net517,net384_c1,dummy52);
wire dummy53;
SPLITT SplitCLK_2_432(net809,net383_c1,dummy53);
wire dummy54;
SPLITT SplitCLK_2_433(net711,net382_c1,dummy54);
wire dummy55;
SPLITT SplitCLK_2_434(net575,net381_c1,dummy55);
wire dummy56;
SPLITT SplitCLK_2_435(net455,net380_c1,dummy56);
wire dummy57;
SPLITT SplitCLK_2_436(net799,net379_c1,dummy57);
wire dummy58;
SPLITT SplitCLK_4_437(net448,net378_c1,dummy58);
wire dummy59;
SPLITT SplitCLK_2_438(net763,net377_c1,dummy59);
wire dummy60;
SPLITT SplitCLK_2_439(net635,net376_c1,dummy60);
wire dummy61;
SPLITT SplitCLK_4_440(net636,net375_c1,dummy61);
wire dummy62;
SPLITT SplitCLK_2_441(net491,net374_c1,dummy62);
wire dummy63;
SPLITT SplitCLK_2_442(net679,net373_c1,dummy63);
wire dummy64;
SPLITT SplitCLK_2_443(net643,net372_c1,dummy64);
wire dummy65;
SPLITT SplitCLK_2_444(net611,net371_c1,dummy65);
SPLITT SplitCLK_0_445(net813,net369_c1,net370_c1);
wire dummy66;
SPLITT Split_HOLD_541(net279,dummy66,net814_c1);
INTERCONNECT DFFT_178_TDO_TDO_Pad(net0_c1,TDO_Pad);
INTERCONNECT TMS_Pad_Split_197_n479(TMS_Pad,net1);
INTERCONNECT NOTT_8_n20_Split_200_n482(net2_c1,net2);
INTERCONNECT AND2T_9_n21_Split_203_n485(net3_c1,net3);
INTERCONNECT AND2T_18_n30_Split_218_n500(net4_c1,net4);
INTERCONNECT NOTT_10_n22_AND2T_96_n114(net5_c1,net5);
INTERCONNECT AND2T_19_n31_DFFT_127__FPB_n409(net6_c1,net6);
INTERCONNECT NOTT_11_n23_Split_205_n487(net7_c1,net7);
INTERCONNECT OR2T_28_n40_OR2T_29_n41(net8_c1,net8);
INTERCONNECT XOR2T_20_n32_AND2T_19_n31(net9_c1,net9);
INTERCONNECT AND2T_12_n24_Split_207_n489(net10_c1,net10);
INTERCONNECT OR2T_29_n41_DFFT_145__FPB_n427(net11_c1,net11);
INTERCONNECT AND2T_21_n33_DFFT_162__FPB_n444(net12_c1,net12);
INTERCONNECT AND2T_13_n25_Split_209_n491(net13_c1,net13);
INTERCONNECT AND2T_38_n50_OR2T_39_n51(net14_c1,net14);
INTERCONNECT AND2T_30_n42_Split_226_n508(net15_c1,net15);
INTERCONNECT AND2T_22_n34_Split_221_n503(net16_c1,net16);
INTERCONNECT AND2T_14_n26_Split_210_n492(net17_c1,net17);
INTERCONNECT OR2T_39_n51_OR2T_50_n62(net18_c1,net18);
INTERCONNECT AND2T_31_n43_Split_229_n511(net19_c1,net19);
INTERCONNECT AND2T_23_n35_Split_222_n504(net20_c1,net20);
INTERCONNECT AND2T_15_n27_Split_213_n495(net21_c1,net21);
INTERCONNECT NOTT_7_n19_AND2T_95_n113(net22_c1,net22);
INTERCONNECT AND2T_48_n60_OR2T_49_n61(net23_c1,net23);
INTERCONNECT AND2T_40_n52_OR2T_42_n54(net24_c1,net24);
INTERCONNECT OR2T_32_n44_AND2T_33_n45(net25_c1,net25);
INTERCONNECT NOTT_24_n36_Split_224_n506(net26_c1,net26);
INTERCONNECT AND2T_16_n28_Split_215_n497(net27_c1,net27);
INTERCONNECT OR2T_49_n61_OR2T_50_n62(net28_c1,net28);
INTERCONNECT AND2T_41_n53_OR2T_42_n54(net29_c1,net29);
INTERCONNECT AND2T_33_n45_OR2T_39_n51(net30_c1,net30);
INTERCONNECT AND2T_25_n37_AND2T_26_n38(net31_c1,net31);
INTERCONNECT AND2T_17_n29_Split_217_n499(net32_c1,net32);
INTERCONNECT AND2T_58_n70_Split_237_n519(net33_c1,net33);
INTERCONNECT OR2T_50_n62_OR2T_51_n63(net34_c1,net34);
INTERCONNECT OR2T_42_n54_Split_233_n515(net35_c1,net35);
INTERCONNECT AND2T_34_n46_Split_230_n512(net36_c1,net36);
INTERCONNECT AND2T_26_n38_Split_225_n507(net37_c1,net37);
INTERCONNECT AND2T_59_n71_Split_238_n520(net38_c1,net38);
INTERCONNECT OR2T_51_n63_DFFT_103__FBL_n385(net39_c1,net39);
INTERCONNECT AND2T_43_n55_OR2T_49_n61(net40_c1,net40);
INTERCONNECT AND2T_35_n47_Split_231_n513(net41_c1,net41);
INTERCONNECT OR2T_27_n39_OR2T_28_n40(net42_c1,net42);
INTERCONNECT OR2T_68_n80_Split_241_n523(net43_c1,net43);
INTERCONNECT OR2T_60_n72_OR2T_66_n78(net44_c1,net44);
INTERCONNECT OR2T_52_n64_Split_236_n518(net45_c1,net45);
INTERCONNECT AND2T_44_n56_Split_234_n516(net46_c1,net46);
INTERCONNECT OR2T_36_n48_AND2T_38_n50(net47_c1,net47);
INTERCONNECT AND2T_69_n81_Split_242_n524(net48_c1,net48);
INTERCONNECT AND2T_61_n73_Split_239_n521(net49_c1,net49);
INTERCONNECT OR2T_53_n65_AND2T_54_n66(net50_c1,net50);
INTERCONNECT AND2T_45_n57_OR2T_47_n59(net51_c1,net51);
INTERCONNECT OR2T_37_n49_AND2T_38_n50(net52_c1,net52);
INTERCONNECT OR2T_78_n90_Split_244_n526(net53_c1,net53);
INTERCONNECT AND2T_70_n82_DFFT_159__FPB_n441(net54_c1,net54);
INTERCONNECT AND2T_62_n74_OR2T_65_n77(net55_c1,net55);
INTERCONNECT AND2T_54_n66_DFFT_157__FPB_n439(net56_c1,net56);
INTERCONNECT AND2T_46_n58_DFFT_141__FPB_n423(net57_c1,net57);
INTERCONNECT AND2T_79_n91_OR2T_82_n94(net58_c1,net58);
INTERCONNECT OR2T_71_n83_OR2T_72_n84(net59_c1,net59);
INTERCONNECT AND2T_63_n75_AND2T_64_n76(net60_c1,net60);
INTERCONNECT AND2T_55_n67_DFFT_150__FPB_n432(net61_c1,net61);
INTERCONNECT OR2T_47_n59_Split_235_n517(net62_c1,net62);
INTERCONNECT OR2T_80_n92_AND2T_79_n91(net63_c1,net63);
INTERCONNECT OR2T_72_n84_DFFT_161__FPB_n443(net64_c1,net64);
INTERCONNECT AND2T_64_n76_Split_240_n522(net65_c1,net65);
INTERCONNECT AND2T_56_n68_AND2T_55_n67(net66_c1,net66);
INTERCONNECT AND2T_81_n93_OR2T_82_n94(net67_c1,net67);
INTERCONNECT OR2T_73_n85_OR2T_77_n89(net68_c1,net68);
INTERCONNECT OR2T_65_n77_OR2T_66_n78(net69_c1,net69);
INTERCONNECT OR2T_57_n69_DFFT_155__FPB_n437(net70_c1,net70);
INTERCONNECT OR2T_82_n94_OR2T_83_n95(net71_c1,net71);
INTERCONNECT AND2T_74_n86_DFFT_160__FPB_n442(net72_c1,net72);
INTERCONNECT OR2T_66_n78_OR2T_67_n79(net73_c1,net73);
INTERCONNECT OR2T_83_n95_DFFT_172__FPB_n454(net74_c1,net74);
INTERCONNECT AND2T_75_n87_AND2T_74_n86(net75_c1,net75);
INTERCONNECT OR2T_67_n79_OR2T_68_n80(net76_c1,net76);
INTERCONNECT AND2T_84_n96_OR2T_86_n98(net77_c1,net77);
INTERCONNECT OR2T_76_n88_OR2T_77_n89(net78_c1,net78);
INTERCONNECT AND2T_85_n97_OR2T_86_n98(net79_c1,net79);
INTERCONNECT OR2T_77_n89_OR2T_78_n90(net80_c1,net80);
INTERCONNECT OR2T_86_n98_OR2T_90_n102(net81_c1,net81);
INTERCONNECT AND2T_87_n99_OR2T_89_n101(net82_c1,net82);
INTERCONNECT AND2T_88_n100_OR2T_89_n101(net83_c1,net83);
INTERCONNECT OR2T_89_n101_OR2T_90_n102(net84_c1,net84);
INTERCONNECT OR2T_90_n102_OR2T_91_n103(net85_c1,net85);
INTERCONNECT OR2T_91_n103_Split_246_n528(net86_c1,net86);
INTERCONNECT AND2T_92_n104_DFFT_179__FPB_n461(net87_c1,net87);
INTERCONNECT AND2T_95_n113_Split_248_n530(net88_c1,net88);
INTERCONNECT AND2T_93_n105_DFFT_185__FPB_n467(net89_c1,net89);
INTERCONNECT AND2T_96_n114_Split_251_n533(net90_c1,net90);
INTERCONNECT AND2T_94_n106_DFFT_191__FPB_n473(net91_c1,net91);
INTERCONNECT NOTT_99_n123_Split_260_n542(net92_c1,net92);
INTERCONNECT AND2T_97_n115_Split_254_n536(net93_c1,net93);
INTERCONNECT NOTT_100_n124_Split_263_n545(net94_c1,net94);
INTERCONNECT NOTT_98_n116_Split_257_n539(net95_c1,net95);
INTERCONNECT Split_218_n500_Split_220_n502(net96_c1,net96);
INTERCONNECT Split_219_n501_AND2T_34_n46(net97_c1,net97);
INTERCONNECT Split_220_n502_AND2T_74_n86(net98_c1,net98);
INTERCONNECT Split_228_n510_AND2T_63_n75(net99_c1,net99);
INTERCONNECT Split_229_n511_OR2T_52_n64(net100_c1,net100);
INTERCONNECT Split_221_n503_OR2T_52_n64(net101_c1,net101);
INTERCONNECT Split_222_n504_Split_223_n505(net102_c1,net102);
INTERCONNECT Split_238_n520_OR2T_76_n88(net103_c1,net103);
INTERCONNECT Split_230_n512_OR2T_71_n83(net104_c1,net104);
INTERCONNECT Split_231_n513_Split_232_n514(net105_c1,net105);
INTERCONNECT Split_239_n521_AND2T_87_n99(net106_c1,net106);
INTERCONNECT Split_223_n505_AND2T_70_n82(net107_c1,net107);
INTERCONNECT Split_248_n530_Split_250_n532(net108_c1,net108);
INTERCONNECT Split_240_n522_OR2T_83_n95(net109_c1,net109);
INTERCONNECT Split_224_n506_DFFT_153__FPB_n435(net110_c1,net110);
INTERCONNECT Split_232_n514_OR2T_37_n49(net111_c1,net111);
INTERCONNECT Split_241_n523_DFFT_107__FBL_n389(net112_c1,net112);
INTERCONNECT Split_233_n515_OR2T_73_n85(net113_c1,net113);
INTERCONNECT Split_225_n507_OR2T_57_n69(net114_c1,net114);
INTERCONNECT Split_249_n531_AND2T_22_n34(net115_c1,net115);
INTERCONNECT Split_226_n508_Split_228_n510(net116_c1,net116);
INTERCONNECT Split_242_n524_Split_243_n525(net117_c1,net117);
INTERCONNECT Split_234_n516_DFFT_154__FPB_n436(net118_c1,net118);
INTERCONNECT Split_250_n532_AND2T_45_n57(net119_c1,net119);
INTERCONNECT Split_258_n540_DFFT_131__FPB_n413(net120_c1,net120);
INTERCONNECT Split_251_n533_Split_253_n535(net121_c1,net121);
INTERCONNECT Split_259_n541_DFFT_151__FPB_n433(net122_c1,net122);
INTERCONNECT Split_243_n525_DFFT_165__FPB_n447(net123_c1,net123);
INTERCONNECT Split_235_n517_OR2T_53_n65(net124_c1,net124);
INTERCONNECT Split_227_n509_AND2T_35_n47(net125_c1,net125);
INTERCONNECT Split_260_n542_Split_262_n544(net126_c1,net126);
INTERCONNECT Split_268_n550_DFFT_137__FPB_n419(net127_c1,net127);
INTERCONNECT Split_244_n526_Split_245_n527(net128_c1,net128);
INTERCONNECT Split_236_n518_OR2T_73_n85(net129_c1,net129);
INTERCONNECT Split_252_n534_AND2T_35_n47(net130_c1,net130);
INTERCONNECT Split_269_n551_Split_271_n553(net131_c1,net131);
INTERCONNECT Split_245_n527_DFFT_116__FPB_n398(net132_c1,net132);
INTERCONNECT Split_237_n519_AND2T_85_n97(net133_c1,net133);
INTERCONNECT Split_253_n535_AND2T_61_n73(net134_c1,net134);
INTERCONNECT Split_261_n543_AND2T_18_n30(net135_c1,net135);
INTERCONNECT Split_254_n536_Split_256_n538(net136_c1,net136);
INTERCONNECT Split_246_n528_Split_247_n529(net137_c1,net137);
INTERCONNECT Split_198_n480_DFFT_101__FPB_n128(net138_c1,net138);
INTERCONNECT Split_270_n552_AND2T_75_n87(net139_c1,net139);
INTERCONNECT Split_262_n544_OR2T_80_n92(net140_c1,net140);
INTERCONNECT Split_278_n560_AND2T_15_n27(net141_c1,net141);
INTERCONNECT Split_263_n545_Split_265_n547(net142_c1,net142);
INTERCONNECT Split_271_n553_DFFT_166__FPB_n448(net143_c1,net143);
INTERCONNECT Split_279_n561_DFFT_125__FPB_n407(net144_c1,net144);
INTERCONNECT Split_247_n529_DFFT_114__FPB_n396(net145_c1,net145);
INTERCONNECT Split_199_n481_DFFT_168__FPB_n450(net146_c1,net146);
INTERCONNECT Split_255_n537_AND2T_75_n87(net147_c1,net147);
INTERCONNECT Split_280_n562_Split_282_n564(net148_c1,net148);
INTERCONNECT Split_272_n554_Split_274_n556(net149_c1,net149);
INTERCONNECT Split_200_n482_Split_202_n484(net150_c1,net150);
INTERCONNECT Split_256_n538_DFFT_130__FPB_n412(net151_c1,net151);
INTERCONNECT Split_208_n490_AND2T_93_n105(net152_c1,net152);
INTERCONNECT Split_264_n546_XOR2T_20_n32(net153_c1,net153);
INTERCONNECT Split_257_n539_Split_259_n541(net154_c1,net154);
INTERCONNECT Split_209_n491_DFFT_173__FPB_n455(net155_c1,net155);
INTERCONNECT Split_265_n547_AND2T_44_n56(net156_c1,net156);
INTERCONNECT Split_281_n563_AND2T_21_n33(net157_c1,net157);
INTERCONNECT Split_201_n483_AND2T_30_n42(net158_c1,net158);
INTERCONNECT Split_273_n555_AND2T_15_n27(net159_c1,net159);
INTERCONNECT Split_266_n548_Split_268_n550(net160_c1,net160);
INTERCONNECT Split_210_n492_Split_212_n494(net161_c1,net161);
INTERCONNECT Split_282_n564_DFFT_126__FPB_n408(net162_c1,net162);
INTERCONNECT Split_274_n556_DFFT_129__FPB_n411(net163_c1,net163);
INTERCONNECT Split_202_n484_AND2T_95_n113(net164_c1,net164);
INTERCONNECT Split_283_n565_Split_285_n567(net165_c1,net165);
INTERCONNECT Split_275_n557_Split_276_n558(net166_c1,net166);
INTERCONNECT Split_203_n485_Split_204_n486(net167_c1,net167);
INTERCONNECT Split_267_n549_DFFT_120__FPB_n402(net168_c1,net168);
INTERCONNECT Split_211_n493_AND2T_34_n46(net169_c1,net169);
INTERCONNECT Split_276_n558_DFFT_158__FPB_n440(net170_c1,net170);
INTERCONNECT Split_204_n486_AND2T_93_n105(net171_c1,net171);
INTERCONNECT Split_212_n494_AND2T_58_n70(net172_c1,net172);
INTERCONNECT Split_284_n566_AND2T_21_n33(net173_c1,net173);
INTERCONNECT Split_277_n559_Split_279_n561(net174_c1,net174);
INTERCONNECT Split_197_n479_Split_199_n481(net175_c1,net175);
INTERCONNECT Split_213_n495_Split_214_n496(net176_c1,net176);
INTERCONNECT Split_205_n487_Split_206_n488(net177_c1,net177);
INTERCONNECT Split_285_n567_DFFT_118__FPB_n400(net178_c1,net178);
INTERCONNECT Split_214_n496_DFFT_119__FPB_n401(net179_c1,net179);
INTERCONNECT Split_206_n488_AND2T_14_n26(net180_c1,net180);
INTERCONNECT Split_207_n489_Split_208_n490(net181_c1,net181);
INTERCONNECT Split_215_n497_Split_216_n498(net182_c1,net182);
INTERCONNECT Split_216_n498_OR2T_71_n83(net183_c1,net183);
INTERCONNECT Split_217_n499_DFFT_128__FPB_n410(net184_c1,net184);
INTERCONNECT Split_218_n500_Split_219_n501(net185_c1,net185);
INTERCONNECT Split_219_n501_AND2T_19_n31(net186_c1,net186);
INTERCONNECT Split_228_n510_AND2T_58_n70(net187_c1,net187);
INTERCONNECT Split_220_n502_AND2T_61_n73(net188_c1,net188);
INTERCONNECT Split_229_n511_OR2T_32_n44(net189_c1,net189);
INTERCONNECT Split_221_n503_OR2T_27_n39(net190_c1,net190);
INTERCONNECT Split_238_n520_OR2T_60_n72(net191_c1,net191);
INTERCONNECT Split_222_n504_AND2T_81_n93(net192_c1,net192);
INTERCONNECT Split_230_n512_OR2T_36_n48(net193_c1,net193);
INTERCONNECT Split_239_n521_AND2T_62_n74(net194_c1,net194);
INTERCONNECT Split_223_n505_AND2T_26_n38(net195_c1,net195);
INTERCONNECT Split_231_n513_AND2T_88_n100(net196_c1,net196);
INTERCONNECT Split_248_n530_Split_249_n531(net197_c1,net197);
INTERCONNECT Split_224_n506_AND2T_63_n75(net198_c1,net198);
INTERCONNECT Split_232_n514_OR2T_36_n48(net199_c1,net199);
INTERCONNECT Split_240_n522_OR2T_65_n77(net200_c1,net200);
INTERCONNECT Split_249_n531_AND2T_13_n25(net201_c1,net201);
INTERCONNECT Split_225_n507_OR2T_27_n39(net202_c1,net202);
INTERCONNECT Split_233_n515_AND2T_43_n55(net203_c1,net203);
INTERCONNECT Split_241_n523_DFFT_104__FBL_n386(net204_c1,net204);
INTERCONNECT Split_258_n540_AND2T_25_n37(net205_c1,net205);
INTERCONNECT Split_226_n508_Split_227_n509(net206_c1,net206);
INTERCONNECT Split_234_n516_AND2T_45_n57(net207_c1,net207);
INTERCONNECT Split_242_n524_DFFT_171__FPB_n453(net208_c1,net208);
INTERCONNECT Split_250_n532_AND2T_41_n53(net209_c1,net209);
INTERCONNECT Split_259_n541_DFFT_142__FPB_n424(net210_c1,net210);
INTERCONNECT Split_227_n509_AND2T_31_n43(net211_c1,net211);
INTERCONNECT Split_235_n517_AND2T_48_n60(net212_c1,net212);
INTERCONNECT Split_243_n525_AND2T_70_n82(net213_c1,net213);
INTERCONNECT Split_251_n533_Split_252_n534(net214_c1,net214);
INTERCONNECT Split_268_n550_DFFT_134__FPB_n416(net215_c1,net215);
INTERCONNECT Split_236_n518_OR2T_53_n65(net216_c1,net216);
INTERCONNECT Split_244_n526_DFFT_117__FPB_n399(net217_c1,net217);
INTERCONNECT Split_252_n534_AND2T_13_n25(net218_c1,net218);
INTERCONNECT Split_260_n542_Split_261_n543(net219_c1,net219);
INTERCONNECT Split_269_n551_Split_270_n552(net220_c1,net220);
INTERCONNECT Split_237_n519_AND2T_59_n71(net221_c1,net221);
INTERCONNECT Split_245_n527_DFFT_112__FPB_n394(net222_c1,net222);
INTERCONNECT Split_253_n535_AND2T_40_n52(net223_c1,net223);
INTERCONNECT Split_261_n543_AND2T_9_n21(net224_c1,net224);
INTERCONNECT Split_198_n480_NOTT_98_n116(net225_c1,net225);
INTERCONNECT Split_278_n560_NOTT_8_n20(net226_c1,net226);
INTERCONNECT Split_246_n528_DFFT_115__FPB_n397(net227_c1,net227);
INTERCONNECT Split_254_n536_Split_255_n537(net228_c1,net228);
INTERCONNECT Split_262_n544_AND2T_55_n67(net229_c1,net229);
INTERCONNECT Split_270_n552_AND2T_69_n81(net230_c1,net230);
INTERCONNECT Split_199_n481_DFFT_102__FPB_n129(net231_c1,net231);
INTERCONNECT Split_279_n561_DFFT_122__FPB_n404(net232_c1,net232);
INTERCONNECT Split_247_n529_DFFT_113__FPB_n395(net233_c1,net233);
INTERCONNECT Split_255_n537_AND2T_46_n58(net234_c1,net234);
INTERCONNECT Split_263_n545_Split_264_n546(net235_c1,net235);
INTERCONNECT Split_271_n553_DFFT_146__FPB_n428(net236_c1,net236);
INTERCONNECT Split_256_n538_DFFT_124__FPB_n406(net237_c1,net237);
INTERCONNECT Split_264_n546_AND2T_12_n24(net238_c1,net238);
INTERCONNECT Split_272_n554_Split_273_n555(net239_c1,net239);
INTERCONNECT Split_280_n562_Split_281_n563(net240_c1,net240);
INTERCONNECT Split_208_n490_AND2T_92_n104(net241_c1,net241);
INTERCONNECT Split_200_n482_Split_201_n483(net242_c1,net242);
INTERCONNECT Split_257_n539_Split_258_n540(net243_c1,net243);
INTERCONNECT Split_265_n547_AND2T_23_n35(net244_c1,net244);
INTERCONNECT Split_273_n555_NOTT_7_n19(net245_c1,net245);
INTERCONNECT Split_281_n563_NOTT_11_n23(net246_c1,net246);
INTERCONNECT Split_209_n491_OR2T_32_n44(net247_c1,net247);
INTERCONNECT Split_201_n483_AND2T_9_n21(net248_c1,net248);
INTERCONNECT Split_266_n548_Split_267_n549(net249_c1,net249);
INTERCONNECT Split_274_n556_NOTT_99_n123(net250_c1,net250);
INTERCONNECT Split_282_n564_DFFT_123__FPB_n405(net251_c1,net251);
INTERCONNECT Split_202_n484_OR2T_80_n92(net252_c1,net252);
INTERCONNECT Split_210_n492_Split_211_n493(net253_c1,net253);
INTERCONNECT Split_267_n549_NOTT_24_n36(net254_c1,net254);
INTERCONNECT Split_275_n557_DFFT_163__FPB_n445(net255_c1,net255);
INTERCONNECT Split_283_n565_Split_284_n566(net256_c1,net256);
INTERCONNECT Split_203_n485_AND2T_94_n106(net257_c1,net257);
INTERCONNECT Split_211_n493_AND2T_16_n28(net258_c1,net258);
INTERCONNECT Split_276_n558_DFFT_140__FPB_n422(net259_c1,net259);
INTERCONNECT Split_284_n566_NOTT_10_n22(net260_c1,net260);
INTERCONNECT Split_204_n486_AND2T_92_n104(net261_c1,net261);
INTERCONNECT Split_212_n494_AND2T_41_n53(net262_c1,net262);
INTERCONNECT Split_197_n479_Split_198_n480(net263_c1,net263);
INTERCONNECT Split_277_n559_Split_278_n560(net264_c1,net264);
INTERCONNECT Split_285_n567_AND2T_56_n68(net265_c1,net265);
INTERCONNECT Split_205_n487_AND2T_96_n114(net266_c1,net266);
INTERCONNECT Split_213_n495_DFFT_136__FPB_n418(net267_c1,net267);
INTERCONNECT Split_206_n488_AND2T_12_n24(net268_c1,net268);
INTERCONNECT Split_214_n496_AND2T_46_n58(net269_c1,net269);
INTERCONNECT Split_207_n489_AND2T_94_n106(net270_c1,net270);
INTERCONNECT Split_215_n497_AND2T_84_n96(net271_c1,net271);
INTERCONNECT Split_216_n498_AND2T_17_n29(net272_c1,net272);
INTERCONNECT Split_217_n499_OR2T_60_n72(net273_c1,net273);
INTERCONNECT DFFT_184_St_obs0_St_obs0_Pad(net274_c1,St_obs0_Pad);
INTERCONNECT DFFT_190_St_obs1_St_obs1_Pad(net275_c1,St_obs1_Pad);
INTERCONNECT DFFT_196_St_obs2_St_obs2_Pad(net276_c1,St_obs2_Pad);
INTERCONNECT DFFT_108__FBL_n390_AND2T_97_n115(net277_c1,net277);
INTERCONNECT DFFT_109__FBL_n391_Split_280_n562(net278_c1,net278);
INTERCONNECT DFFT_110__FBL_n392_Split_HOLD_541(net279_c1,net279);
INTERCONNECT DFFT_111__FBL_n393_Split_283_n565(net280_c1,net280);
INTERCONNECT DFFT_103__FBL_n385_Split_272_n554(net281_c1,net281);
INTERCONNECT DFFT_104__FBL_n386_AND2T_56_n68(net282_c1,net282);
INTERCONNECT DFFT_105__FBL_n387_AND2T_97_n115(net283_c1,net283);
INTERCONNECT DFFT_106__FBL_n388_Split_275_n557(net284_c1,net284);
INTERCONNECT DFFT_107__FBL_n389_Split_277_n559(net285_c1,net285);
INTERCONNECT DFFT_101__FPB_n128_Split_266_n548(net286_c1,net286);
INTERCONNECT DFFT_118__FPB_n400_AND2T_14_n26(net287_c1,net287);
INTERCONNECT DFFT_102__FPB_n129_Split_269_n551(net288_c1,net288);
INTERCONNECT DFFT_119__FPB_n401_AND2T_16_n28(net289_c1,net289);
INTERCONNECT DFFT_120__FPB_n402_DFFT_121__FPB_n403(net290_c1,net290);
INTERCONNECT DFFT_128__FPB_n410_OR2T_29_n41(net291_c1,net291);
INTERCONNECT DFFT_129__FPB_n411_AND2T_30_n42(net292_c1,net292);
INTERCONNECT DFFT_121__FPB_n403_AND2T_17_n29(net293_c1,net293);
INTERCONNECT DFFT_138__FPB_n420_DFFT_139__FPB_n421(net294_c1,net294);
INTERCONNECT DFFT_130__FPB_n412_AND2T_31_n43(net295_c1,net295);
INTERCONNECT DFFT_122__FPB_n404_AND2T_18_n30(net296_c1,net296);
INTERCONNECT DFFT_131__FPB_n413_DFFT_132__FPB_n414(net297_c1,net297);
INTERCONNECT DFFT_139__FPB_n421_AND2T_43_n55(net298_c1,net298);
INTERCONNECT DFFT_123__FPB_n405_XOR2T_20_n32(net299_c1,net299);
INTERCONNECT DFFT_148__FPB_n430_DFFT_149__FPB_n431(net300_c1,net300);
INTERCONNECT DFFT_132__FPB_n414_DFFT_133__FPB_n415(net301_c1,net301);
INTERCONNECT DFFT_140__FPB_n422_AND2T_44_n56(net302_c1,net302);
INTERCONNECT DFFT_124__FPB_n406_AND2T_22_n34(net303_c1,net303);
INTERCONNECT DFFT_149__FPB_n431_AND2T_54_n66(net304_c1,net304);
INTERCONNECT DFFT_141__FPB_n423_OR2T_47_n59(net305_c1,net305);
INTERCONNECT DFFT_133__FPB_n415_AND2T_33_n45(net306_c1,net306);
INTERCONNECT DFFT_125__FPB_n407_AND2T_23_n35(net307_c1,net307);
INTERCONNECT DFFT_142__FPB_n424_DFFT_143__FPB_n425(net308_c1,net308);
INTERCONNECT DFFT_134__FPB_n416_DFFT_135__FPB_n417(net309_c1,net309);
INTERCONNECT DFFT_158__FPB_n440_AND2T_69_n81(net310_c1,net310);
INTERCONNECT DFFT_150__FPB_n432_OR2T_57_n69(net311_c1,net311);
INTERCONNECT DFFT_126__FPB_n408_AND2T_25_n37(net312_c1,net312);
INTERCONNECT DFFT_151__FPB_n433_DFFT_152__FPB_n434(net313_c1,net313);
INTERCONNECT DFFT_143__FPB_n425_DFFT_144__FPB_n426(net314_c1,net314);
INTERCONNECT DFFT_159__FPB_n441_OR2T_72_n84(net315_c1,net315);
INTERCONNECT DFFT_135__FPB_n417_OR2T_37_n49(net316_c1,net316);
INTERCONNECT DFFT_127__FPB_n409_OR2T_28_n40(net317_c1,net317);
INTERCONNECT DFFT_168__FPB_n450_DFFT_169__FPB_n451(net318_c1,net318);
INTERCONNECT DFFT_160__FPB_n442_OR2T_76_n88(net319_c1,net319);
INTERCONNECT DFFT_152__FPB_n434_AND2T_59_n71(net320_c1,net320);
INTERCONNECT DFFT_144__FPB_n426_AND2T_48_n60(net321_c1,net321);
INTERCONNECT DFFT_136__FPB_n418_AND2T_40_n52(net322_c1,net322);
INTERCONNECT DFFT_169__FPB_n451_DFFT_170__FPB_n452(net323_c1,net323);
INTERCONNECT DFFT_137__FPB_n419_DFFT_138__FPB_n420(net324_c1,net324);
INTERCONNECT DFFT_161__FPB_n443_OR2T_78_n90(net325_c1,net325);
INTERCONNECT DFFT_153__FPB_n435_AND2T_62_n74(net326_c1,net326);
INTERCONNECT DFFT_145__FPB_n427_OR2T_51_n63(net327_c1,net327);
INTERCONNECT DFFT_146__FPB_n428_DFFT_147__FPB_n429(net328_c1,net328);
INTERCONNECT DFFT_170__FPB_n452_AND2T_87_n99(net329_c1,net329);
INTERCONNECT DFFT_162__FPB_n444_AND2T_79_n91(net330_c1,net330);
INTERCONNECT DFFT_154__FPB_n436_AND2T_64_n76(net331_c1,net331);
INTERCONNECT DFFT_179__FPB_n461_DFFT_180__FPB_n462(net332_c1,net332);
INTERCONNECT DFFT_163__FPB_n445_DFFT_164__FPB_n446(net333_c1,net333);
INTERCONNECT DFFT_155__FPB_n437_DFFT_156__FPB_n438(net334_c1,net334);
INTERCONNECT DFFT_147__FPB_n429_DFFT_148__FPB_n430(net335_c1,net335);
INTERCONNECT DFFT_171__FPB_n453_AND2T_88_n100(net336_c1,net336);
INTERCONNECT DFFT_188__FPB_n470_DFFT_189__FPB_n471(net337_c1,net337);
INTERCONNECT DFFT_180__FPB_n462_DFFT_181__FPB_n463(net338_c1,net338);
INTERCONNECT DFFT_172__FPB_n454_OR2T_91_n103(net339_c1,net339);
INTERCONNECT DFFT_164__FPB_n446_AND2T_81_n93(net340_c1,net340);
INTERCONNECT DFFT_156__FPB_n438_OR2T_67_n79(net341_c1,net341);
INTERCONNECT DFFT_189__FPB_n471_DFFT_190_St_obs1(net342_c1,net342);
INTERCONNECT DFFT_181__FPB_n463_DFFT_182__FPB_n464(net343_c1,net343);
INTERCONNECT DFFT_173__FPB_n455_DFFT_174__FPB_n456(net344_c1,net344);
INTERCONNECT DFFT_165__FPB_n447_AND2T_84_n96(net345_c1,net345);
INTERCONNECT DFFT_157__FPB_n439_OR2T_68_n80(net346_c1,net346);
INTERCONNECT DFFT_182__FPB_n464_DFFT_183__FPB_n465(net347_c1,net347);
INTERCONNECT DFFT_174__FPB_n456_DFFT_175__FPB_n457(net348_c1,net348);
INTERCONNECT DFFT_166__FPB_n448_DFFT_167__FPB_n449(net349_c1,net349);
INTERCONNECT DFFT_191__FPB_n473_DFFT_192__FPB_n474(net350_c1,net350);
INTERCONNECT DFFT_183__FPB_n465_DFFT_184_St_obs0(net351_c1,net351);
INTERCONNECT DFFT_175__FPB_n457_DFFT_176__FPB_n458(net352_c1,net352);
INTERCONNECT DFFT_167__FPB_n449_AND2T_85_n97(net353_c1,net353);
INTERCONNECT DFFT_192__FPB_n474_DFFT_193__FPB_n475(net354_c1,net354);
INTERCONNECT DFFT_176__FPB_n458_DFFT_177__FPB_n459(net355_c1,net355);
INTERCONNECT DFFT_112__FPB_n394_DFFT_105__FBL_n387(net356_c1,net356);
INTERCONNECT DFFT_193__FPB_n475_DFFT_194__FPB_n476(net357_c1,net357);
INTERCONNECT DFFT_185__FPB_n467_DFFT_186__FPB_n468(net358_c1,net358);
INTERCONNECT DFFT_177__FPB_n459_DFFT_178_TDO(net359_c1,net359);
INTERCONNECT DFFT_113__FPB_n395_DFFT_106__FBL_n388(net360_c1,net360);
INTERCONNECT DFFT_194__FPB_n476_DFFT_195__FPB_n477(net361_c1,net361);
INTERCONNECT DFFT_186__FPB_n468_DFFT_187__FPB_n469(net362_c1,net362);
INTERCONNECT DFFT_114__FPB_n396_DFFT_108__FBL_n390(net363_c1,net363);
INTERCONNECT DFFT_195__FPB_n477_DFFT_196_St_obs2(net364_c1,net364);
INTERCONNECT DFFT_187__FPB_n469_DFFT_188__FPB_n470(net365_c1,net365);
INTERCONNECT DFFT_115__FPB_n397_DFFT_109__FBL_n391(net366_c1,net366);
INTERCONNECT DFFT_116__FPB_n398_DFFT_110__FBL_n392(net367_c1,net367);
INTERCONNECT DFFT_117__FPB_n399_DFFT_111__FBL_n393(net368_c1,net368);
INTERCONNECT SplitCLK_0_445_SplitCLK_0_284(net369_c1,net369);
INTERCONNECT SplitCLK_0_445_SplitCLK_2_378(net370_c1,net370);
INTERCONNECT SplitCLK_2_444_NOTT_98_n116(net371_c1,net371);
INTERCONNECT SplitCLK_2_443_DFFT_187__FPB_n469(net372_c1,net372);
INTERCONNECT SplitCLK_2_442_DFFT_195__FPB_n477(net373_c1,net373);
INTERCONNECT SplitCLK_2_441_DFFT_179__FPB_n461(net374_c1,net374);
INTERCONNECT SplitCLK_4_440_DFFT_186__FPB_n468(net375_c1,net375);
INTERCONNECT SplitCLK_2_439_DFFT_185__FPB_n467(net376_c1,net376);
INTERCONNECT SplitCLK_2_438_DFFT_169__FPB_n451(net377_c1,net377);
INTERCONNECT SplitCLK_4_437_DFFT_183__FPB_n465(net378_c1,net378);
INTERCONNECT SplitCLK_2_436_DFFT_166__FPB_n448(net379_c1,net379);
INTERCONNECT SplitCLK_2_435_DFFT_182__FPB_n464(net380_c1,net380);
INTERCONNECT SplitCLK_2_434_DFFT_173__FPB_n455(net381_c1,net381);
INTERCONNECT SplitCLK_2_433_DFFT_164__FPB_n446(net382_c1,net382);
INTERCONNECT SplitCLK_2_432_DFFT_147__FPB_n429(net383_c1,net383);
INTERCONNECT SplitCLK_2_431_DFFT_155__FPB_n437(net384_c1,net384);
INTERCONNECT SplitCLK_2_430_DFFT_154__FPB_n436(net385_c1,net385);
INTERCONNECT SplitCLK_2_429_DFFT_137__FPB_n419(net386_c1,net386);
INTERCONNECT SplitCLK_2_428_DFFT_153__FPB_n435(net387_c1,net387);
INTERCONNECT SplitCLK_2_427_DFFT_161__FPB_n443(net388_c1,net388);
INTERCONNECT SplitCLK_2_426_DFFT_136__FPB_n418(net389_c1,net389);
INTERCONNECT SplitCLK_2_425_DFFT_128__FPB_n410(net390_c1,net390);
INTERCONNECT SplitCLK_2_424_DFFT_127__FPB_n409(net391_c1,net391);
INTERCONNECT SplitCLK_2_423_DFFT_135__FPB_n417(net392_c1,net392);
INTERCONNECT SplitCLK_2_422_DFFT_143__FPB_n425(net393_c1,net393);
INTERCONNECT SplitCLK_2_421_DFFT_142__FPB_n424(net394_c1,net394);
INTERCONNECT SplitCLK_2_420_DFFT_125__FPB_n407(net395_c1,net395);
INTERCONNECT SplitCLK_2_419_DFFT_133__FPB_n415(net396_c1,net396);
INTERCONNECT SplitCLK_4_418_DFFT_108__FBL_n390(net397_c1,net397);
INTERCONNECT SplitCLK_2_417_DFFT_115__FPB_n397(net398_c1,net398);
INTERCONNECT SplitCLK_2_416_DFFT_107__FBL_n389(net399_c1,net399);
INTERCONNECT SplitCLK_4_415_DFFT_105__FBL_n387(net400_c1,net400);
INTERCONNECT SplitCLK_2_414_DFFT_112__FPB_n394(net401_c1,net401);
INTERCONNECT SplitCLK_2_413_DFFT_120__FPB_n402(net402_c1,net402);
INTERCONNECT SplitCLK_2_412_DFFT_111__FBL_n393(net403_c1,net403);
INTERCONNECT SplitCLK_2_411_DFFT_110__FBL_n392(net404_c1,net404);
INTERCONNECT SplitCLK_2_410_AND2T_96_n114(net405_c1,net405);
INTERCONNECT SplitCLK_2_409_AND2T_95_n113(net406_c1,net406);
INTERCONNECT SplitCLK_2_408_AND2T_92_n104(net407_c1,net407);
INTERCONNECT SplitCLK_2_407_NOTT_24_n36(net408_c1,net408);
INTERCONNECT SplitCLK_2_406_OR2T_67_n79(net409_c1,net409);
INTERCONNECT SplitCLK_2_405_DFFT_178_TDO(net410_c1,net410);
INTERCONNECT SplitCLK_2_404_OR2T_66_n78(net411_c1,net411);
INTERCONNECT SplitCLK_2_403_OR2T_49_n61(net412_c1,net412);
INTERCONNECT SplitCLK_2_402_OR2T_72_n84(net413_c1,net413);
INTERCONNECT SplitCLK_2_401_OR2T_80_n92(net414_c1,net414);
INTERCONNECT SplitCLK_2_400_OR2T_39_n51(net415_c1,net415);
INTERCONNECT SplitCLK_2_399_OR2T_29_n41(net416_c1,net416);
INTERCONNECT SplitCLK_2_398_OR2T_52_n64(net417_c1,net417);
INTERCONNECT SplitCLK_2_397_OR2T_51_n63(net418_c1,net418);
INTERCONNECT SplitCLK_2_396_OR2T_42_n54(net419_c1,net419);
INTERCONNECT SplitCLK_4_395_AND2T_85_n97(net420_c1,net420);
INTERCONNECT SplitCLK_2_394_AND2T_74_n86(net421_c1,net421);
INTERCONNECT SplitCLK_2_393_AND2T_56_n68(net422_c1,net422);
INTERCONNECT SplitCLK_4_392_AND2T_64_n76(net423_c1,net423);
INTERCONNECT SplitCLK_4_391_AND2T_46_n58(net424_c1,net424);
INTERCONNECT SplitCLK_2_390_AND2T_54_n66(net425_c1,net425);
INTERCONNECT SplitCLK_2_389_AND2T_43_n55(net426_c1,net426);
INTERCONNECT SplitCLK_2_388_AND2T_19_n31(net427_c1,net427);
INTERCONNECT SplitCLK_2_387_AND2T_26_n38(net428_c1,net428);
INTERCONNECT SplitCLK_2_386_AND2T_34_n46(net429_c1,net429);
INTERCONNECT SplitCLK_2_385_AND2T_17_n29(net430_c1,net430);
INTERCONNECT SplitCLK_2_384_AND2T_14_n26(net431_c1,net431);
INTERCONNECT SplitCLK_4_383_AND2T_22_n34(net432_c1,net432);
INTERCONNECT SplitCLK_2_382_AND2T_13_n25(net433_c1,net433);
INTERCONNECT SplitCLK_2_381_AND2T_21_n33(net434_c1,net434);
INTERCONNECT SplitCLK_2_380_DFFT_184_St_obs0(net435_c1,net435);
INTERCONNECT SplitCLK_2_379_AND2T_9_n21(net436_c1,net436);
INTERCONNECT SplitCLK_2_378_SplitCLK_6_331(net437_c1,net437);
INTERCONNECT SplitCLK_2_378_SplitCLK_4_377(net438_c1,net438);
INTERCONNECT SplitCLK_4_377_SplitCLK_0_354(net439_c1,net439);
INTERCONNECT SplitCLK_4_377_SplitCLK_2_376(net440_c1,net440);
INTERCONNECT SplitCLK_2_376_SplitCLK_6_365(net441_c1,net441);
INTERCONNECT SplitCLK_2_376_SplitCLK_4_375(net442_c1,net442);
INTERCONNECT SplitCLK_4_375_SplitCLK_0_370(net443_c1,net443);
INTERCONNECT SplitCLK_4_375_SplitCLK_2_374(net444_c1,net444);
INTERCONNECT SplitCLK_2_374_SplitCLK_6_372(net445_c1,net445);
INTERCONNECT SplitCLK_2_374_SplitCLK_4_373(net446_c1,net446);
INTERCONNECT SplitCLK_4_373_SplitCLK_2_380(net447_c1,net447);
INTERCONNECT SplitCLK_4_373_SplitCLK_4_437(net448_c1,net448);
INTERCONNECT SplitCLK_6_372_SplitCLK_2_410(net449_c1,net449);
INTERCONNECT SplitCLK_6_372_SplitCLK_4_371(net450_c1,net450);
INTERCONNECT SplitCLK_4_371_NOTT_10_n22(net451_c1,net451);
INTERCONNECT SplitCLK_4_371_NOTT_11_n23(net452_c1,net452);
INTERCONNECT SplitCLK_0_370_SplitCLK_6_367(net453_c1,net453);
INTERCONNECT SplitCLK_0_370_SplitCLK_4_369(net454_c1,net454);
INTERCONNECT SplitCLK_4_369_SplitCLK_2_435(net455_c1,net455);
INTERCONNECT SplitCLK_4_369_SplitCLK_4_368(net456_c1,net456);
INTERCONNECT SplitCLK_4_368_DFFT_180__FPB_n462(net457_c1,net457);
INTERCONNECT SplitCLK_4_368_DFFT_181__FPB_n463(net458_c1,net458);
INTERCONNECT SplitCLK_6_367_SplitCLK_2_381(net459_c1,net459);
INTERCONNECT SplitCLK_6_367_SplitCLK_4_366(net460_c1,net460);
INTERCONNECT SplitCLK_4_366_AND2T_79_n91(net461_c1,net461);
INTERCONNECT SplitCLK_4_366_DFFT_162__FPB_n444(net462_c1,net462);
INTERCONNECT SplitCLK_6_365_SplitCLK_0_359(net463_c1,net463);
INTERCONNECT SplitCLK_6_365_SplitCLK_4_364(net464_c1,net464);
INTERCONNECT SplitCLK_4_364_SplitCLK_2_361(net465_c1,net465);
INTERCONNECT SplitCLK_4_364_SplitCLK_4_363(net466_c1,net466);
INTERCONNECT SplitCLK_4_363_SplitCLK_2_409(net467_c1,net467);
INTERCONNECT SplitCLK_4_363_SplitCLK_4_362(net468_c1,net468);
INTERCONNECT SplitCLK_4_362_NOTT_7_n19(net469_c1,net469);
INTERCONNECT SplitCLK_4_362_NOTT_8_n20(net470_c1,net470);
INTERCONNECT SplitCLK_2_361_SplitCLK_2_426(net471_c1,net471);
INTERCONNECT SplitCLK_2_361_SplitCLK_4_360(net472_c1,net472);
INTERCONNECT SplitCLK_4_360_DFFT_103__FBL_n385(net473_c1,net473);
INTERCONNECT SplitCLK_4_360_DFFT_129__FPB_n411(net474_c1,net474);
INTERCONNECT SplitCLK_0_359_SplitCLK_2_356(net475_c1,net475);
INTERCONNECT SplitCLK_0_359_SplitCLK_2_358(net476_c1,net476);
INTERCONNECT SplitCLK_2_358_SplitCLK_2_401(net477_c1,net477);
INTERCONNECT SplitCLK_2_358_SplitCLK_4_357(net478_c1,net478);
INTERCONNECT SplitCLK_4_357_AND2T_30_n42(net479_c1,net479);
INTERCONNECT SplitCLK_4_357_NOTT_99_n123(net480_c1,net480);
INTERCONNECT SplitCLK_2_356_SplitCLK_2_396(net481_c1,net481);
INTERCONNECT SplitCLK_2_356_SplitCLK_4_355(net482_c1,net482);
INTERCONNECT SplitCLK_4_355_OR2T_27_n39(net483_c1,net483);
INTERCONNECT SplitCLK_4_355_OR2T_57_n69(net484_c1,net484);
INTERCONNECT SplitCLK_0_354_SplitCLK_6_342(net485_c1,net485);
INTERCONNECT SplitCLK_0_354_SplitCLK_4_353(net486_c1,net486);
INTERCONNECT SplitCLK_4_353_SplitCLK_0_347(net487_c1,net487);
INTERCONNECT SplitCLK_4_353_SplitCLK_2_352(net488_c1,net488);
INTERCONNECT SplitCLK_2_352_SplitCLK_2_349(net489_c1,net489);
INTERCONNECT SplitCLK_2_352_SplitCLK_4_351(net490_c1,net490);
INTERCONNECT SplitCLK_4_351_SplitCLK_2_441(net491_c1,net491);
INTERCONNECT SplitCLK_4_351_SplitCLK_4_350(net492_c1,net492);
INTERCONNECT SplitCLK_4_350_DFFT_190_St_obs1(net493_c1,net493);
INTERCONNECT SplitCLK_4_350_DFFT_189__FPB_n471(net494_c1,net494);
INTERCONNECT SplitCLK_2_349_SplitCLK_2_384(net495_c1,net495);
INTERCONNECT SplitCLK_2_349_SplitCLK_4_348(net496_c1,net496);
INTERCONNECT SplitCLK_4_348_AND2T_12_n24(net497_c1,net497);
INTERCONNECT SplitCLK_4_348_DFFT_118__FPB_n400(net498_c1,net498);
INTERCONNECT SplitCLK_0_347_SplitCLK_6_344(net499_c1,net499);
INTERCONNECT SplitCLK_0_347_SplitCLK_2_346(net500_c1,net500);
INTERCONNECT SplitCLK_2_346_SplitCLK_2_408(net501_c1,net501);
INTERCONNECT SplitCLK_2_346_SplitCLK_4_345(net502_c1,net502);
INTERCONNECT SplitCLK_4_345_AND2T_93_n105(net503_c1,net503);
INTERCONNECT SplitCLK_4_345_AND2T_94_n106(net504_c1,net504);
INTERCONNECT SplitCLK_6_344_SplitCLK_2_393(net505_c1,net505);
INTERCONNECT SplitCLK_6_344_SplitCLK_4_343(net506_c1,net506);
INTERCONNECT SplitCLK_4_343_XOR2T_20_n32(net507_c1,net507);
INTERCONNECT SplitCLK_4_343_DFFT_123__FPB_n405(net508_c1,net508);
INTERCONNECT SplitCLK_6_342_SplitCLK_0_336(net509_c1,net509);
INTERCONNECT SplitCLK_6_342_SplitCLK_6_341(net510_c1,net510);
INTERCONNECT SplitCLK_6_341_SplitCLK_4_338(net511_c1,net511);
INTERCONNECT SplitCLK_6_341_SplitCLK_4_340(net512_c1,net512);
INTERCONNECT SplitCLK_4_340_SplitCLK_2_424(net513_c1,net513);
INTERCONNECT SplitCLK_4_340_SplitCLK_4_339(net514_c1,net514);
INTERCONNECT SplitCLK_4_339_AND2T_15_n27(net515_c1,net515);
INTERCONNECT SplitCLK_4_339_AND2T_55_n67(net516_c1,net516);
INTERCONNECT SplitCLK_4_338_SplitCLK_2_431(net517_c1,net517);
INTERCONNECT SplitCLK_4_338_SplitCLK_4_337(net518_c1,net518);
INTERCONNECT SplitCLK_4_337_AND2T_41_n53(net519_c1,net519);
INTERCONNECT SplitCLK_4_337_DFFT_156__FPB_n438(net520_c1,net520);
INTERCONNECT SplitCLK_0_336_SplitCLK_6_333(net521_c1,net521);
INTERCONNECT SplitCLK_0_336_SplitCLK_2_335(net522_c1,net522);
INTERCONNECT SplitCLK_2_335_SplitCLK_2_379(net523_c1,net523);
INTERCONNECT SplitCLK_2_335_SplitCLK_4_334(net524_c1,net524);
INTERCONNECT SplitCLK_4_334_DFFT_104__FBL_n386(net525_c1,net525);
INTERCONNECT SplitCLK_4_334_DFFT_150__FPB_n432(net526_c1,net526);
INTERCONNECT SplitCLK_6_333_SplitCLK_2_406(net527_c1,net527);
INTERCONNECT SplitCLK_6_333_SplitCLK_4_332(net528_c1,net528);
INTERCONNECT SplitCLK_4_332_AND2T_45_n57(net529_c1,net529);
INTERCONNECT SplitCLK_4_332_OR2T_68_n80(net530_c1,net530);
INTERCONNECT SplitCLK_6_331_SplitCLK_0_307(net531_c1,net531);
INTERCONNECT SplitCLK_6_331_SplitCLK_6_330(net532_c1,net532);
INTERCONNECT SplitCLK_6_330_SplitCLK_6_318(net533_c1,net533);
INTERCONNECT SplitCLK_6_330_SplitCLK_4_329(net534_c1,net534);
INTERCONNECT SplitCLK_4_329_SplitCLK_0_323(net535_c1,net535);
INTERCONNECT SplitCLK_4_329_SplitCLK_4_328(net536_c1,net536);
INTERCONNECT SplitCLK_4_328_SplitCLK_2_325(net537_c1,net537);
INTERCONNECT SplitCLK_4_328_SplitCLK_4_327(net538_c1,net538);
INTERCONNECT SplitCLK_4_327_SplitCLK_2_382(net539_c1,net539);
INTERCONNECT SplitCLK_4_327_SplitCLK_4_326(net540_c1,net540);
INTERCONNECT SplitCLK_4_326_AND2T_40_n52(net541_c1,net541);
INTERCONNECT SplitCLK_4_326_DFFT_124__FPB_n406(net542_c1,net542);
INTERCONNECT SplitCLK_2_325_SplitCLK_2_398(net543_c1,net543);
INTERCONNECT SplitCLK_2_325_SplitCLK_4_324(net544_c1,net544);
INTERCONNECT SplitCLK_4_324_OR2T_37_n49(net545_c1,net545);
INTERCONNECT SplitCLK_4_324_DFFT_130__FPB_n412(net546_c1,net546);
INTERCONNECT SplitCLK_0_323_SplitCLK_2_320(net547_c1,net547);
INTERCONNECT SplitCLK_0_323_SplitCLK_4_322(net548_c1,net548);
INTERCONNECT SplitCLK_4_322_SplitCLK_4_383(net549_c1,net549);
INTERCONNECT SplitCLK_4_322_SplitCLK_4_321(net550_c1,net550);
INTERCONNECT SplitCLK_4_321_AND2T_31_n43(net551_c1,net551);
INTERCONNECT SplitCLK_4_321_AND2T_35_n47(net552_c1,net552);
INTERCONNECT SplitCLK_2_320_SplitCLK_2_389(net553_c1,net553);
INTERCONNECT SplitCLK_2_320_SplitCLK_4_319(net554_c1,net554);
INTERCONNECT SplitCLK_4_319_AND2T_38_n50(net555_c1,net555);
INTERCONNECT SplitCLK_4_319_OR2T_73_n85(net556_c1,net556);
INTERCONNECT SplitCLK_6_318_SplitCLK_4_312(net557_c1,net557);
INTERCONNECT SplitCLK_6_318_SplitCLK_6_317(net558_c1,net558);
INTERCONNECT SplitCLK_6_317_SplitCLK_6_314(net559_c1,net559);
INTERCONNECT SplitCLK_6_317_SplitCLK_2_316(net560_c1,net560);
INTERCONNECT SplitCLK_2_316_SplitCLK_2_423(net561_c1,net561);
INTERCONNECT SplitCLK_2_316_SplitCLK_4_315(net562_c1,net562);
INTERCONNECT SplitCLK_4_315_OR2T_32_n44(net563_c1,net563);
INTERCONNECT SplitCLK_4_315_DFFT_134__FPB_n416(net564_c1,net564);
INTERCONNECT SplitCLK_6_314_SplitCLK_2_405(net565_c1,net565);
INTERCONNECT SplitCLK_6_314_SplitCLK_4_313(net566_c1,net566);
INTERCONNECT SplitCLK_4_313_DFFT_176__FPB_n458(net567_c1,net567);
INTERCONNECT SplitCLK_4_313_DFFT_177__FPB_n459(net568_c1,net568);
INTERCONNECT SplitCLK_4_312_SplitCLK_6_309(net569_c1,net569);
INTERCONNECT SplitCLK_4_312_SplitCLK_6_311(net570_c1,net570);
INTERCONNECT SplitCLK_6_311_SplitCLK_2_429(net571_c1,net571);
INTERCONNECT SplitCLK_6_311_SplitCLK_4_310(net572_c1,net572);
INTERCONNECT SplitCLK_4_310_DFFT_138__FPB_n420(net573_c1,net573);
INTERCONNECT SplitCLK_4_310_DFFT_139__FPB_n421(net574_c1,net574);
INTERCONNECT SplitCLK_6_309_SplitCLK_2_434(net575_c1,net575);
INTERCONNECT SplitCLK_6_309_SplitCLK_4_308(net576_c1,net576);
INTERCONNECT SplitCLK_4_308_DFFT_174__FPB_n456(net577_c1,net577);
INTERCONNECT SplitCLK_4_308_DFFT_175__FPB_n457(net578_c1,net578);
INTERCONNECT SplitCLK_0_307_SplitCLK_6_295(net579_c1,net579);
INTERCONNECT SplitCLK_0_307_SplitCLK_4_306(net580_c1,net580);
INTERCONNECT SplitCLK_4_306_SplitCLK_0_300(net581_c1,net581);
INTERCONNECT SplitCLK_4_306_SplitCLK_6_305(net582_c1,net582);
INTERCONNECT SplitCLK_6_305_SplitCLK_6_302(net583_c1,net583);
INTERCONNECT SplitCLK_6_305_SplitCLK_2_304(net584_c1,net584);
INTERCONNECT SplitCLK_2_304_SplitCLK_2_399(net585_c1,net585);
INTERCONNECT SplitCLK_2_304_SplitCLK_4_303(net586_c1,net586);
INTERCONNECT SplitCLK_4_303_AND2T_58_n70(net587_c1,net587);
INTERCONNECT SplitCLK_4_303_OR2T_28_n40(net588_c1,net588);
INTERCONNECT SplitCLK_6_302_SplitCLK_2_397(net589_c1,net589);
INTERCONNECT SplitCLK_6_302_SplitCLK_4_301(net590_c1,net590);
INTERCONNECT SplitCLK_4_301_AND2T_59_n71(net591_c1,net591);
INTERCONNECT SplitCLK_4_301_DFFT_145__FPB_n427(net592_c1,net592);
INTERCONNECT SplitCLK_0_300_SplitCLK_6_297(net593_c1,net593);
INTERCONNECT SplitCLK_0_300_SplitCLK_4_299(net594_c1,net594);
INTERCONNECT SplitCLK_4_299_SplitCLK_2_404(net595_c1,net595);
INTERCONNECT SplitCLK_4_299_SplitCLK_4_298(net596_c1,net596);
INTERCONNECT SplitCLK_4_298_AND2T_61_n73(net597_c1,net597);
INTERCONNECT SplitCLK_4_298_DFFT_160__FPB_n442(net598_c1,net598);
INTERCONNECT SplitCLK_6_297_SplitCLK_2_425(net599_c1,net599);
INTERCONNECT SplitCLK_6_297_SplitCLK_4_296(net600_c1,net600);
INTERCONNECT SplitCLK_4_296_OR2T_60_n72(net601_c1,net601);
INTERCONNECT SplitCLK_4_296_OR2T_77_n89(net602_c1,net602);
INTERCONNECT SplitCLK_6_295_SplitCLK_0_289(net603_c1,net603);
INTERCONNECT SplitCLK_6_295_SplitCLK_6_294(net604_c1,net604);
INTERCONNECT SplitCLK_6_294_SplitCLK_6_291(net605_c1,net605);
INTERCONNECT SplitCLK_6_294_SplitCLK_4_293(net606_c1,net606);
INTERCONNECT SplitCLK_4_293_SplitCLK_2_419(net607_c1,net607);
INTERCONNECT SplitCLK_4_293_SplitCLK_4_292(net608_c1,net608);
INTERCONNECT SplitCLK_4_292_AND2T_33_n45(net609_c1,net609);
INTERCONNECT SplitCLK_4_292_OR2T_36_n48(net610_c1,net610);
INTERCONNECT SplitCLK_6_291_SplitCLK_2_444(net611_c1,net611);
INTERCONNECT SplitCLK_6_291_SplitCLK_4_290(net612_c1,net612);
INTERCONNECT SplitCLK_4_290_DFFT_131__FPB_n413(net613_c1,net613);
INTERCONNECT SplitCLK_4_290_DFFT_132__FPB_n414(net614_c1,net614);
INTERCONNECT SplitCLK_0_289_SplitCLK_4_286(net615_c1,net615);
INTERCONNECT SplitCLK_0_289_SplitCLK_2_288(net616_c1,net616);
INTERCONNECT SplitCLK_2_288_SplitCLK_2_400(net617_c1,net617);
INTERCONNECT SplitCLK_2_288_SplitCLK_4_287(net618_c1,net618);
INTERCONNECT SplitCLK_4_287_OR2T_50_n62(net619_c1,net619);
INTERCONNECT SplitCLK_4_287_DFFT_157__FPB_n439(net620_c1,net620);
INTERCONNECT SplitCLK_4_286_SplitCLK_2_422(net621_c1,net621);
INTERCONNECT SplitCLK_4_286_SplitCLK_4_285(net622_c1,net622);
INTERCONNECT SplitCLK_4_285_DFFT_101__FPB_n128(net623_c1,net623);
INTERCONNECT SplitCLK_4_285_DFFT_144__FPB_n426(net624_c1,net624);
INTERCONNECT SplitCLK_0_284_SplitCLK_6_237(net625_c1,net625);
INTERCONNECT SplitCLK_0_284_SplitCLK_4_283(net626_c1,net626);
INTERCONNECT SplitCLK_4_283_SplitCLK_0_260(net627_c1,net627);
INTERCONNECT SplitCLK_4_283_SplitCLK_2_282(net628_c1,net628);
INTERCONNECT SplitCLK_2_282_SplitCLK_2_271(net629_c1,net629);
INTERCONNECT SplitCLK_2_282_SplitCLK_4_281(net630_c1,net630);
INTERCONNECT SplitCLK_4_281_SplitCLK_0_276(net631_c1,net631);
INTERCONNECT SplitCLK_4_281_SplitCLK_6_280(net632_c1,net632);
INTERCONNECT SplitCLK_6_280_SplitCLK_4_278(net633_c1,net633);
INTERCONNECT SplitCLK_6_280_SplitCLK_4_279(net634_c1,net634);
INTERCONNECT SplitCLK_4_279_SplitCLK_2_439(net635_c1,net635);
INTERCONNECT SplitCLK_4_279_SplitCLK_4_440(net636_c1,net636);
INTERCONNECT SplitCLK_4_278_SplitCLK_2_412(net637_c1,net637);
INTERCONNECT SplitCLK_4_278_SplitCLK_4_277(net638_c1,net638);
INTERCONNECT SplitCLK_4_277_DFFT_109__FBL_n391(net639_c1,net639);
INTERCONNECT SplitCLK_4_277_DFFT_117__FPB_n399(net640_c1,net640);
INTERCONNECT SplitCLK_0_276_SplitCLK_2_273(net641_c1,net641);
INTERCONNECT SplitCLK_0_276_SplitCLK_4_275(net642_c1,net642);
INTERCONNECT SplitCLK_4_275_SplitCLK_2_443(net643_c1,net643);
INTERCONNECT SplitCLK_4_275_SplitCLK_4_274(net644_c1,net644);
INTERCONNECT SplitCLK_4_274_DFFT_196_St_obs2(net645_c1,net645);
INTERCONNECT SplitCLK_4_274_DFFT_188__FPB_n470(net646_c1,net646);
INTERCONNECT SplitCLK_2_273_SplitCLK_2_417(net647_c1,net647);
INTERCONNECT SplitCLK_2_273_SplitCLK_4_272(net648_c1,net648);
INTERCONNECT SplitCLK_4_272_AND2T_97_n115(net649_c1,net649);
INTERCONNECT SplitCLK_4_272_NOTT_100_n124(net650_c1,net650);
INTERCONNECT SplitCLK_2_271_SplitCLK_4_265(net651_c1,net651);
INTERCONNECT SplitCLK_2_271_SplitCLK_2_270(net652_c1,net652);
INTERCONNECT SplitCLK_2_270_SplitCLK_2_267(net653_c1,net653);
INTERCONNECT SplitCLK_2_270_SplitCLK_4_269(net654_c1,net654);
INTERCONNECT SplitCLK_4_269_SplitCLK_2_416(net655_c1,net655);
INTERCONNECT SplitCLK_4_269_SplitCLK_4_268(net656_c1,net656);
INTERCONNECT SplitCLK_4_268_DFFT_122__FPB_n404(net657_c1,net657);
INTERCONNECT SplitCLK_4_268_DFFT_126__FPB_n408(net658_c1,net658);
INTERCONNECT SplitCLK_2_267_SplitCLK_2_388(net659_c1,net659);
INTERCONNECT SplitCLK_2_267_SplitCLK_4_266(net660_c1,net660);
INTERCONNECT SplitCLK_4_266_AND2T_25_n37(net661_c1,net661);
INTERCONNECT SplitCLK_4_266_OR2T_47_n59(net662_c1,net662);
INTERCONNECT SplitCLK_4_265_SplitCLK_4_262(net663_c1,net663);
INTERCONNECT SplitCLK_4_265_SplitCLK_2_264(net664_c1,net664);
INTERCONNECT SplitCLK_2_264_SplitCLK_2_420(net665_c1,net665);
INTERCONNECT SplitCLK_2_264_SplitCLK_4_263(net666_c1,net666);
INTERCONNECT SplitCLK_4_263_AND2T_23_n35(net667_c1,net667);
INTERCONNECT SplitCLK_4_263_AND2T_18_n30(net668_c1,net668);
INTERCONNECT SplitCLK_4_262_SplitCLK_2_387(net669_c1,net669);
INTERCONNECT SplitCLK_4_262_SplitCLK_4_261(net670_c1,net670);
INTERCONNECT SplitCLK_4_261_AND2T_16_n28(net671_c1,net671);
INTERCONNECT SplitCLK_4_261_AND2T_44_n56(net672_c1,net672);
INTERCONNECT SplitCLK_0_260_SplitCLK_6_248(net673_c1,net673);
INTERCONNECT SplitCLK_0_260_SplitCLK_4_259(net674_c1,net674);
INTERCONNECT SplitCLK_4_259_SplitCLK_4_253(net675_c1,net675);
INTERCONNECT SplitCLK_4_259_SplitCLK_2_258(net676_c1,net676);
INTERCONNECT SplitCLK_2_258_SplitCLK_6_255(net677_c1,net677);
INTERCONNECT SplitCLK_2_258_SplitCLK_4_257(net678_c1,net678);
INTERCONNECT SplitCLK_4_257_SplitCLK_2_442(net679_c1,net679);
INTERCONNECT SplitCLK_4_257_SplitCLK_4_256(net680_c1,net680);
INTERCONNECT SplitCLK_4_256_DFFT_193__FPB_n475(net681_c1,net681);
INTERCONNECT SplitCLK_4_256_DFFT_194__FPB_n476(net682_c1,net682);
INTERCONNECT SplitCLK_6_255_SplitCLK_2_411(net683_c1,net683);
INTERCONNECT SplitCLK_6_255_SplitCLK_4_254(net684_c1,net684);
INTERCONNECT SplitCLK_4_254_DFFT_114__FPB_n396(net685_c1,net685);
INTERCONNECT SplitCLK_4_254_DFFT_116__FPB_n398(net686_c1,net686);
INTERCONNECT SplitCLK_4_253_SplitCLK_0_250(net687_c1,net687);
INTERCONNECT SplitCLK_4_253_SplitCLK_4_252(net688_c1,net688);
INTERCONNECT SplitCLK_4_252_SplitCLK_2_414(net689_c1,net689);
INTERCONNECT SplitCLK_4_252_SplitCLK_4_251(net690_c1,net690);
INTERCONNECT SplitCLK_4_251_DFFT_191__FPB_n473(net691_c1,net691);
INTERCONNECT SplitCLK_4_251_DFFT_192__FPB_n474(net692_c1,net692);
INTERCONNECT SplitCLK_0_250_SplitCLK_4_415(net693_c1,net693);
INTERCONNECT SplitCLK_0_250_SplitCLK_4_249(net694_c1,net694);
INTERCONNECT SplitCLK_4_249_DFFT_113__FPB_n395(net695_c1,net695);
INTERCONNECT SplitCLK_4_249_DFFT_106__FBL_n388(net696_c1,net696);
INTERCONNECT SplitCLK_6_248_SplitCLK_0_242(net697_c1,net697);
INTERCONNECT SplitCLK_6_248_SplitCLK_2_247(net698_c1,net698);
INTERCONNECT SplitCLK_2_247_SplitCLK_6_244(net699_c1,net699);
INTERCONNECT SplitCLK_2_247_SplitCLK_4_246(net700_c1,net700);
INTERCONNECT SplitCLK_4_246_SplitCLK_4_418(net701_c1,net701);
INTERCONNECT SplitCLK_4_246_SplitCLK_4_245(net702_c1,net702);
INTERCONNECT SplitCLK_4_245_AND2T_81_n93(net703_c1,net703);
INTERCONNECT SplitCLK_4_245_OR2T_82_n94(net704_c1,net704);
INTERCONNECT SplitCLK_6_244_SplitCLK_2_386(net705_c1,net705);
INTERCONNECT SplitCLK_6_244_SplitCLK_4_243(net706_c1,net706);
INTERCONNECT SplitCLK_4_243_OR2T_83_n95(net707_c1,net707);
INTERCONNECT SplitCLK_4_243_DFFT_172__FPB_n454(net708_c1,net708);
INTERCONNECT SplitCLK_0_242_SplitCLK_6_239(net709_c1,net709);
INTERCONNECT SplitCLK_0_242_SplitCLK_2_241(net710_c1,net710);
INTERCONNECT SplitCLK_2_241_SplitCLK_2_433(net711_c1,net711);
INTERCONNECT SplitCLK_2_241_SplitCLK_4_240(net712_c1,net712);
INTERCONNECT SplitCLK_4_240_OR2T_91_n103(net713_c1,net713);
INTERCONNECT SplitCLK_4_240_DFFT_163__FPB_n445(net714_c1,net714);
INTERCONNECT SplitCLK_6_239_SplitCLK_2_430(net715_c1,net715);
INTERCONNECT SplitCLK_6_239_SplitCLK_4_238(net716_c1,net716);
INTERCONNECT SplitCLK_4_238_DFFT_140__FPB_n422(net717_c1,net717);
INTERCONNECT SplitCLK_4_238_DFFT_158__FPB_n440(net718_c1,net718);
INTERCONNECT SplitCLK_6_237_SplitCLK_0_213(net719_c1,net719);
INTERCONNECT SplitCLK_6_237_SplitCLK_2_236(net720_c1,net720);
INTERCONNECT SplitCLK_2_236_SplitCLK_6_224(net721_c1,net721);
INTERCONNECT SplitCLK_2_236_SplitCLK_4_235(net722_c1,net722);
INTERCONNECT SplitCLK_4_235_SplitCLK_4_229(net723_c1,net723);
INTERCONNECT SplitCLK_4_235_SplitCLK_2_234(net724_c1,net724);
INTERCONNECT SplitCLK_2_234_SplitCLK_2_231(net725_c1,net725);
INTERCONNECT SplitCLK_2_234_SplitCLK_4_233(net726_c1,net726);
INTERCONNECT SplitCLK_4_233_SplitCLK_2_394(net727_c1,net727);
INTERCONNECT SplitCLK_4_233_SplitCLK_4_232(net728_c1,net728);
INTERCONNECT SplitCLK_4_232_OR2T_78_n90(net729_c1,net729);
INTERCONNECT SplitCLK_4_232_DFFT_141__FPB_n423(net730_c1,net730);
INTERCONNECT SplitCLK_2_231_SplitCLK_2_385(net731_c1,net731);
INTERCONNECT SplitCLK_2_231_SplitCLK_4_230(net732_c1,net732);
INTERCONNECT SplitCLK_4_230_OR2T_71_n83(net733_c1,net733);
INTERCONNECT SplitCLK_4_230_OR2T_76_n88(net734_c1,net734);
INTERCONNECT SplitCLK_4_229_SplitCLK_2_226(net735_c1,net735);
INTERCONNECT SplitCLK_4_229_SplitCLK_2_228(net736_c1,net736);
INTERCONNECT SplitCLK_2_228_SplitCLK_2_427(net737_c1,net737);
INTERCONNECT SplitCLK_2_228_SplitCLK_4_227(net738_c1,net738);
INTERCONNECT SplitCLK_4_227_AND2T_75_n87(net739_c1,net739);
INTERCONNECT SplitCLK_4_227_DFFT_119__FPB_n401(net740_c1,net740);
INTERCONNECT SplitCLK_2_226_SplitCLK_2_402(net741_c1,net741);
INTERCONNECT SplitCLK_2_226_SplitCLK_4_225(net742_c1,net742);
INTERCONNECT SplitCLK_4_225_OR2T_86_n98(net743_c1,net743);
INTERCONNECT SplitCLK_4_225_DFFT_165__FPB_n447(net744_c1,net744);
INTERCONNECT SplitCLK_6_224_SplitCLK_0_218(net745_c1,net745);
INTERCONNECT SplitCLK_6_224_SplitCLK_2_223(net746_c1,net746);
INTERCONNECT SplitCLK_2_223_SplitCLK_2_220(net747_c1,net747);
INTERCONNECT SplitCLK_2_223_SplitCLK_4_222(net748_c1,net748);
INTERCONNECT SplitCLK_4_222_SplitCLK_2_403(net749_c1,net749);
INTERCONNECT SplitCLK_4_222_SplitCLK_4_221(net750_c1,net750);
INTERCONNECT SplitCLK_4_221_AND2T_48_n60(net751_c1,net751);
INTERCONNECT SplitCLK_4_221_AND2T_84_n96(net752_c1,net752);
INTERCONNECT SplitCLK_2_220_SplitCLK_2_421(net753_c1,net753);
INTERCONNECT SplitCLK_2_220_SplitCLK_0_219(net754_c1,net754);
INTERCONNECT SplitCLK_0_219_DFFT_102__FPB_n129(net755_c1,net755);
INTERCONNECT SplitCLK_0_219_DFFT_168__FPB_n450(net756_c1,net756);
INTERCONNECT SplitCLK_0_218_SplitCLK_2_215(net757_c1,net757);
INTERCONNECT SplitCLK_0_218_SplitCLK_4_217(net758_c1,net758);
INTERCONNECT SplitCLK_4_217_SplitCLK_4_395(net759_c1,net759);
INTERCONNECT SplitCLK_4_217_SplitCLK_4_216(net760_c1,net760);
INTERCONNECT SplitCLK_4_216_OR2T_53_n65(net761_c1,net761);
INTERCONNECT SplitCLK_4_216_DFFT_152__FPB_n434(net762_c1,net762);
INTERCONNECT SplitCLK_2_215_SplitCLK_2_438(net763_c1,net763);
INTERCONNECT SplitCLK_2_215_SplitCLK_4_214(net764_c1,net764);
INTERCONNECT SplitCLK_4_214_DFFT_151__FPB_n433(net765_c1,net765);
INTERCONNECT SplitCLK_4_214_DFFT_170__FPB_n452(net766_c1,net766);
INTERCONNECT SplitCLK_0_213_SplitCLK_6_201(net767_c1,net767);
INTERCONNECT SplitCLK_0_213_SplitCLK_4_212(net768_c1,net768);
INTERCONNECT SplitCLK_4_212_SplitCLK_0_206(net769_c1,net769);
INTERCONNECT SplitCLK_4_212_SplitCLK_4_211(net770_c1,net770);
INTERCONNECT SplitCLK_4_211_SplitCLK_6_208(net771_c1,net771);
INTERCONNECT SplitCLK_4_211_SplitCLK_6_210(net772_c1,net772);
INTERCONNECT SplitCLK_6_210_SplitCLK_4_391(net773_c1,net773);
INTERCONNECT SplitCLK_6_210_SplitCLK_4_209(net774_c1,net774);
INTERCONNECT SplitCLK_4_209_AND2T_70_n82(net775_c1,net775);
INTERCONNECT SplitCLK_4_209_DFFT_159__FPB_n441(net776_c1,net776);
INTERCONNECT SplitCLK_6_208_SplitCLK_2_428(net777_c1,net777);
INTERCONNECT SplitCLK_6_208_SplitCLK_4_207(net778_c1,net778);
INTERCONNECT SplitCLK_4_207_AND2T_62_n74(net779_c1,net779);
INTERCONNECT SplitCLK_4_207_AND2T_63_n75(net780_c1,net780);
INTERCONNECT SplitCLK_0_206_SplitCLK_6_203(net781_c1,net781);
INTERCONNECT SplitCLK_0_206_SplitCLK_4_205(net782_c1,net782);
INTERCONNECT SplitCLK_4_205_SplitCLK_4_392(net783_c1,net783);
INTERCONNECT SplitCLK_4_205_SplitCLK_4_204(net784_c1,net784);
INTERCONNECT SplitCLK_4_204_AND2T_69_n81(net785_c1,net785);
INTERCONNECT SplitCLK_4_204_OR2T_65_n77(net786_c1,net786);
INTERCONNECT SplitCLK_6_203_SplitCLK_2_407(net787_c1,net787);
INTERCONNECT SplitCLK_6_203_SplitCLK_4_202(net788_c1,net788);
INTERCONNECT SplitCLK_4_202_AND2T_87_n99(net789_c1,net789);
INTERCONNECT SplitCLK_4_202_DFFT_171__FPB_n453(net790_c1,net790);
INTERCONNECT SplitCLK_6_201_SplitCLK_4_195(net791_c1,net791);
INTERCONNECT SplitCLK_6_201_SplitCLK_6_200(net792_c1,net792);
INTERCONNECT SplitCLK_6_200_SplitCLK_6_197(net793_c1,net793);
INTERCONNECT SplitCLK_6_200_SplitCLK_2_199(net794_c1,net794);
INTERCONNECT SplitCLK_2_199_SplitCLK_2_390(net795_c1,net795);
INTERCONNECT SplitCLK_2_199_SplitCLK_4_198(net796_c1,net796);
INTERCONNECT SplitCLK_4_198_AND2T_88_n100(net797_c1,net797);
INTERCONNECT SplitCLK_4_198_OR2T_90_n102(net798_c1,net798);
INTERCONNECT SplitCLK_6_197_SplitCLK_2_436(net799_c1,net799);
INTERCONNECT SplitCLK_6_197_SplitCLK_4_196(net800_c1,net800);
INTERCONNECT SplitCLK_4_196_DFFT_121__FPB_n403(net801_c1,net801);
INTERCONNECT SplitCLK_4_196_DFFT_146__FPB_n428(net802_c1,net802);
INTERCONNECT SplitCLK_4_195_SplitCLK_0_192(net803_c1,net803);
INTERCONNECT SplitCLK_4_195_SplitCLK_2_194(net804_c1,net804);
INTERCONNECT SplitCLK_2_194_SplitCLK_2_413(net805_c1,net805);
INTERCONNECT SplitCLK_2_194_SplitCLK_4_193(net806_c1,net806);
INTERCONNECT SplitCLK_4_193_OR2T_89_n101(net807_c1,net807);
INTERCONNECT SplitCLK_4_193_DFFT_167__FPB_n449(net808_c1,net808);
INTERCONNECT SplitCLK_0_192_SplitCLK_2_432(net809_c1,net809);
INTERCONNECT SplitCLK_0_192_SplitCLK_4_191(net810_c1,net810);
INTERCONNECT SplitCLK_4_191_DFFT_148__FPB_n430(net811_c1,net811);
INTERCONNECT SplitCLK_4_191_DFFT_149__FPB_n431(net812_c1,net812);
INTERCONNECT GCLK_Pad_SplitCLK_0_445(GCLK_Pad,net813);
INTERCONNECT Split_HOLD_541_NOTT_100_n124(net814_c1,net814);

endmodule
