module TAP_route(
input GCLK_Pad,
input TMS_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output state_obs2_Pad,
output state_obs3_Pad);

wire TMS_Pad;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire TRST_Pad;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire net486_c1;
wire net486;
wire net487_c1;
wire net487;
wire net488_c1;
wire net488;
wire net489_c1;
wire net489;
wire net490_c1;
wire net490;
wire net491_c1;
wire net491;
wire net492_c1;
wire net492;
wire net493_c1;
wire net493;
wire net494_c1;
wire net494;
wire net495_c1;
wire net495;
wire net496_c1;
wire net496;
wire net497_c1;
wire net497;
wire net498_c1;
wire net498;
wire net499_c1;
wire net499;
wire net500_c1;
wire net500;
wire net501_c1;
wire net501;
wire net502_c1;
wire net502;
wire net503_c1;
wire net503;
wire net504_c1;
wire net504;
wire net505_c1;
wire net505;
wire net506_c1;
wire net506;
wire net507_c1;
wire net507;
wire net508_c1;
wire net508;
wire net509_c1;
wire net509;
wire net510_c1;
wire net510;
wire net511_c1;
wire net511;
wire net512_c1;
wire net512;
wire net513_c1;
wire net513;
wire net514_c1;
wire net514;
wire net515_c1;
wire net515;
wire net516_c1;
wire net516;
wire net517_c1;
wire net517;
wire net518_c1;
wire net518;
wire net519_c1;
wire net519;
wire net520_c1;
wire net520;
wire net521_c1;
wire net521;
wire net522_c1;
wire net522;
wire net523_c1;
wire net523;
wire net524_c1;
wire net524;
wire net525_c1;
wire net525;
wire net526_c1;
wire net526;
wire net527_c1;
wire net527;
wire net528_c1;
wire net528;
wire net529_c1;
wire net529;
wire net530_c1;
wire net530;
wire net531_c1;
wire net531;
wire net532_c1;
wire net532;
wire net533_c1;
wire net533;
wire net534_c1;
wire net534;
wire net535_c1;
wire net535;
wire net536_c1;
wire net536;
wire net537_c1;
wire net537;
wire net538_c1;
wire net538;
wire net539_c1;
wire net539;
wire net540_c1;
wire net540;
wire net541_c1;
wire net541;
wire net542_c1;
wire net542;
wire net543_c1;
wire net543;
wire net544_c1;
wire net544;
wire net545_c1;
wire net545;
wire net546_c1;
wire net546;
wire net547_c1;
wire state_obs0_Pad;
wire net548_c1;
wire state_obs1_Pad;
wire net549_c1;
wire state_obs2_Pad;
wire net550_c1;
wire state_obs3_Pad;
wire net551_c1;
wire net551;
wire net552_c1;
wire net552;
wire net553_c1;
wire net553;
wire net554_c1;
wire net554;
wire net555_c1;
wire net555;
wire net556_c1;
wire net556;
wire net557_c1;
wire net557;
wire net558_c1;
wire net558;
wire net559_c1;
wire net559;
wire net560_c1;
wire net560;
wire net561_c1;
wire net561;
wire net562_c1;
wire net562;
wire net563_c1;
wire net563;
wire net564_c1;
wire net564;
wire net565_c1;
wire net565;
wire net566_c1;
wire net566;
wire net567_c1;
wire net567;
wire net568_c1;
wire net568;
wire net569_c1;
wire net569;
wire net570_c1;
wire net570;
wire net571_c1;
wire net571;
wire net572_c1;
wire net572;
wire net573_c1;
wire net573;
wire net574_c1;
wire net574;
wire net575_c1;
wire net575;
wire net576_c1;
wire net576;
wire net577_c1;
wire net577;
wire net578_c1;
wire net578;
wire net579_c1;
wire net579;
wire net580_c1;
wire net580;
wire net581_c1;
wire net581;
wire net582_c1;
wire net582;
wire net583_c1;
wire net583;
wire net584_c1;
wire net584;
wire net585_c1;
wire net585;
wire net586_c1;
wire net586;
wire net587_c1;
wire net587;
wire net588_c1;
wire net588;
wire net589_c1;
wire net589;
wire net590_c1;
wire net590;
wire net591_c1;
wire net591;
wire net592_c1;
wire net592;
wire net593_c1;
wire net593;
wire net594_c1;
wire net594;
wire net595_c1;
wire net595;
wire net596_c1;
wire net596;
wire net597_c1;
wire net597;
wire net598_c1;
wire net598;
wire net599_c1;
wire net599;
wire net600_c1;
wire net600;
wire net601_c1;
wire net601;
wire net602_c1;
wire net602;
wire net603_c1;
wire net603;
wire net604_c1;
wire net604;
wire net605_c1;
wire net605;
wire net606_c1;
wire net606;
wire net607_c1;
wire net607;
wire net608_c1;
wire net608;
wire net609_c1;
wire net609;
wire net610_c1;
wire net610;
wire net611_c1;
wire net611;
wire net612_c1;
wire net612;
wire net613_c1;
wire net613;
wire net614_c1;
wire net614;
wire net615_c1;
wire net615;
wire net616_c1;
wire net616;
wire net617_c1;
wire net617;
wire net618_c1;
wire net618;
wire net619_c1;
wire net619;
wire net620_c1;
wire net620;
wire net621_c1;
wire net621;
wire net622_c1;
wire net622;
wire net623_c1;
wire net623;
wire net624_c1;
wire net624;
wire net625_c1;
wire net625;
wire net626_c1;
wire net626;
wire net627_c1;
wire net627;
wire net628_c1;
wire net628;
wire net629_c1;
wire net629;
wire net630_c1;
wire net630;
wire net631_c1;
wire net631;
wire net632_c1;
wire net632;
wire net633_c1;
wire net633;
wire net634_c1;
wire net634;
wire net635_c1;
wire net635;
wire net636_c1;
wire net636;
wire net637_c1;
wire net637;
wire net638_c1;
wire net638;
wire net639_c1;
wire net639;
wire net640_c1;
wire net640;
wire net641_c1;
wire net641;
wire net642_c1;
wire net642;
wire net643_c1;
wire net643;
wire net644_c1;
wire net644;
wire net645_c1;
wire net645;
wire net646_c1;
wire net646;
wire net647_c1;
wire net647;
wire net648_c1;
wire net648;
wire net649_c1;
wire net649;
wire net650_c1;
wire net650;
wire net651_c1;
wire net651;
wire net652_c1;
wire net652;
wire net653_c1;
wire net653;
wire net654_c1;
wire net654;
wire net655_c1;
wire net655;
wire net656_c1;
wire net656;
wire net657_c1;
wire net657;
wire net658_c1;
wire net658;
wire net659_c1;
wire net659;
wire net660_c1;
wire net660;
wire net661_c1;
wire net661;
wire net662_c1;
wire net662;
wire net663_c1;
wire net663;
wire net664_c1;
wire net664;
wire net665_c1;
wire net665;
wire net666_c1;
wire net666;
wire net667_c1;
wire net667;
wire net668_c1;
wire net668;
wire net669_c1;
wire net669;
wire net670_c1;
wire net670;
wire net671_c1;
wire net671;
wire net672_c1;
wire net672;
wire net673_c1;
wire net673;
wire net674_c1;
wire net674;
wire net675_c1;
wire net675;
wire net676_c1;
wire net676;
wire net677_c1;
wire net677;
wire net678_c1;
wire net678;
wire net679_c1;
wire net679;
wire net680_c1;
wire net680;
wire net681_c1;
wire net681;
wire net682_c1;
wire net682;
wire net683_c1;
wire net683;
wire net684_c1;
wire net684;
wire net685_c1;
wire net685;
wire net686_c1;
wire net686;
wire net687_c1;
wire net687;
wire net688_c1;
wire net688;
wire net689_c1;
wire net689;
wire net690_c1;
wire net690;
wire net691_c1;
wire net691;
wire net692_c1;
wire net692;
wire net693_c1;
wire net693;
wire net694_c1;
wire net694;
wire net695_c1;
wire net695;
wire net696_c1;
wire net696;
wire net697_c1;
wire net697;
wire net698_c1;
wire net698;
wire net699_c1;
wire net699;
wire net700_c1;
wire net700;
wire net701_c1;
wire net701;
wire net702_c1;
wire net702;
wire net703_c1;
wire net703;
wire net704_c1;
wire net704;
wire net705_c1;
wire net705;
wire net706_c1;
wire net706;
wire net707_c1;
wire net707;
wire net708_c1;
wire net708;
wire net709_c1;
wire net709;
wire net710_c1;
wire net710;
wire net711_c1;
wire net711;
wire net712_c1;
wire net712;
wire net713_c1;
wire net713;
wire net714_c1;
wire net714;
wire net715_c1;
wire net715;
wire net716_c1;
wire net716;
wire net717_c1;
wire net717;
wire net718_c1;
wire net718;
wire net719_c1;
wire net719;
wire net720_c1;
wire net720;
wire net721_c1;
wire net721;
wire net722_c1;
wire net722;
wire net723_c1;
wire net723;
wire net724_c1;
wire net724;
wire net725_c1;
wire net725;
wire net726_c1;
wire net726;
wire net727_c1;
wire net727;
wire net728_c1;
wire net728;
wire net729_c1;
wire net729;
wire net730_c1;
wire net730;
wire net731_c1;
wire net731;
wire net732_c1;
wire net732;
wire net733_c1;
wire net733;
wire net734_c1;
wire net734;
wire net735_c1;
wire net735;
wire net736_c1;
wire net736;
wire net737_c1;
wire net737;
wire net738_c1;
wire net738;
wire net739_c1;
wire net739;
wire net740_c1;
wire net740;
wire net741_c1;
wire net741;
wire net742_c1;
wire net742;
wire net743_c1;
wire net743;
wire net744_c1;
wire net744;
wire net745_c1;
wire net745;
wire net746_c1;
wire net746;
wire net747_c1;
wire net747;
wire net748_c1;
wire net748;
wire net749_c1;
wire net749;
wire net750_c1;
wire net750;
wire net751_c1;
wire net751;
wire net752_c1;
wire net752;
wire net753_c1;
wire net753;
wire net754_c1;
wire net754;
wire net755_c1;
wire net755;
wire net756_c1;
wire net756;
wire net757_c1;
wire net757;
wire net758_c1;
wire net758;
wire net759_c1;
wire net759;
wire net760_c1;
wire net760;
wire net761_c1;
wire net761;
wire net762_c1;
wire net762;
wire net763_c1;
wire net763;
wire net764_c1;
wire net764;
wire net765_c1;
wire net765;
wire net766_c1;
wire net766;
wire net767_c1;
wire net767;
wire net768_c1;
wire net768;
wire net769_c1;
wire net769;
wire net770_c1;
wire net770;
wire net771_c1;
wire net771;
wire net772_c1;
wire net772;
wire net773_c1;
wire net773;
wire net774_c1;
wire net774;
wire net775_c1;
wire net775;
wire net776_c1;
wire net776;
wire net777_c1;
wire net777;
wire net778_c1;
wire net778;
wire net779_c1;
wire net779;
wire net780_c1;
wire net780;
wire net781_c1;
wire net781;
wire net782_c1;
wire net782;
wire net783_c1;
wire net783;
wire net784_c1;
wire net784;
wire net785_c1;
wire net785;
wire net786_c1;
wire net786;
wire net787_c1;
wire net787;
wire net788_c1;
wire net788;
wire net789_c1;
wire net789;
wire net790_c1;
wire net790;
wire net791_c1;
wire net791;
wire net792_c1;
wire net792;
wire net793_c1;
wire net793;
wire net794_c1;
wire net794;
wire net795_c1;
wire net795;
wire net796_c1;
wire net796;
wire net797_c1;
wire net797;
wire net798_c1;
wire net798;
wire net799_c1;
wire net799;
wire net800_c1;
wire net800;
wire net801_c1;
wire net801;
wire net802_c1;
wire net802;
wire net803_c1;
wire net803;
wire net804_c1;
wire net804;
wire net805_c1;
wire net805;
wire net806_c1;
wire net806;
wire net807_c1;
wire net807;
wire net808_c1;
wire net808;
wire net809_c1;
wire net809;
wire net810_c1;
wire net810;
wire net811_c1;
wire net811;
wire net812_c1;
wire net812;
wire net813_c1;
wire net813;
wire net814_c1;
wire net814;
wire net815_c1;
wire net815;
wire net816_c1;
wire net816;
wire net817_c1;
wire net817;
wire net818_c1;
wire net818;
wire net819_c1;
wire net819;
wire net820_c1;
wire net820;
wire net821_c1;
wire net821;
wire net822_c1;
wire net822;
wire net823_c1;
wire net823;
wire net824_c1;
wire net824;
wire net825_c1;
wire net825;
wire net826_c1;
wire net826;
wire net827_c1;
wire net827;
wire net828_c1;
wire net828;
wire net829_c1;
wire net829;
wire net830_c1;
wire net830;
wire net831_c1;
wire net831;
wire net832_c1;
wire net832;
wire net833_c1;
wire net833;
wire net834_c1;
wire net834;
wire net835_c1;
wire net835;
wire net836_c1;
wire net836;
wire net837_c1;
wire net837;
wire net838_c1;
wire net838;
wire net839_c1;
wire net839;
wire net840_c1;
wire net840;
wire net841_c1;
wire net841;
wire net842_c1;
wire net842;
wire net843_c1;
wire net843;
wire net844_c1;
wire net844;
wire net845_c1;
wire net845;
wire net846_c1;
wire net846;
wire net847_c1;
wire net847;
wire net848_c1;
wire net848;
wire net849_c1;
wire net849;
wire net850_c1;
wire net850;
wire net851_c1;
wire net851;
wire net852_c1;
wire net852;
wire net853_c1;
wire net853;
wire net854_c1;
wire net854;
wire net855_c1;
wire net855;
wire net856_c1;
wire net856;
wire net857_c1;
wire net857;
wire net858_c1;
wire net858;
wire net859_c1;
wire net859;
wire net860_c1;
wire net860;
wire net861_c1;
wire net861;
wire net862_c1;
wire net862;
wire net863_c1;
wire net863;
wire net864_c1;
wire net864;
wire net865_c1;
wire net865;
wire net866_c1;
wire net866;
wire net867_c1;
wire net867;
wire net868_c1;
wire net868;
wire net869_c1;
wire net869;
wire net870_c1;
wire net870;
wire net871_c1;
wire net871;
wire net872_c1;
wire net872;
wire net873_c1;
wire net873;
wire net874_c1;
wire net874;
wire net875_c1;
wire net875;
wire net876_c1;
wire net876;
wire net877_c1;
wire net877;
wire net878_c1;
wire net878;
wire net879_c1;
wire net879;
wire net880_c1;
wire net880;
wire net881_c1;
wire net881;
wire net882_c1;
wire net882;
wire net883_c1;
wire net883;
wire net884_c1;
wire net884;
wire net885_c1;
wire net885;
wire net886_c1;
wire net886;
wire net887_c1;
wire net887;
wire net888_c1;
wire net888;
wire net889_c1;
wire net889;
wire net890_c1;
wire net890;
wire net891_c1;
wire net891;
wire net892_c1;
wire net892;
wire net893_c1;
wire net893;
wire net894_c1;
wire net894;
wire net895_c1;
wire net895;
wire net896_c1;
wire net896;
wire net897_c1;
wire net897;
wire net898_c1;
wire net898;
wire net899_c1;
wire net899;
wire net900_c1;
wire net900;
wire net901_c1;
wire net901;
wire net902_c1;
wire net902;
wire net903_c1;
wire net903;
wire net904_c1;
wire net904;
wire net905_c1;
wire net905;
wire net906_c1;
wire net906;
wire net907_c1;
wire net907;
wire net908_c1;
wire net908;
wire net909_c1;
wire net909;
wire net910_c1;
wire net910;
wire net911_c1;
wire net911;
wire net912_c1;
wire net912;
wire net913_c1;
wire net913;
wire net914_c1;
wire net914;
wire net915_c1;
wire net915;
wire net916_c1;
wire net916;
wire net917_c1;
wire net917;
wire net918_c1;
wire net918;
wire net919_c1;
wire net919;
wire net920_c1;
wire net920;
wire net921_c1;
wire net921;
wire net922_c1;
wire net922;
wire net923_c1;
wire net923;
wire net924_c1;
wire net924;
wire net925_c1;
wire net925;
wire net926_c1;
wire net926;
wire net927_c1;
wire net927;
wire net928_c1;
wire net928;
wire net929_c1;
wire net929;
wire net930_c1;
wire net930;
wire net931_c1;
wire net931;
wire net932_c1;
wire net932;
wire net933_c1;
wire net933;
wire net934_c1;
wire net934;
wire net935_c1;
wire net935;
wire net936_c1;
wire net936;
wire net937_c1;
wire net937;
wire net938_c1;
wire net938;
wire net939_c1;
wire net939;
wire net940_c1;
wire net940;
wire net941_c1;
wire net941;
wire net942_c1;
wire net942;
wire net943_c1;
wire net943;
wire net944_c1;
wire net944;
wire net945_c1;
wire net945;
wire net946_c1;
wire net946;
wire net947_c1;
wire net947;
wire net948_c1;
wire net948;
wire net949_c1;
wire net949;
wire net950_c1;
wire net950;
wire net951_c1;
wire net951;
wire net952_c1;
wire net952;
wire net953_c1;
wire net953;
wire net954_c1;
wire net954;
wire net955_c1;
wire net955;
wire net956_c1;
wire net956;
wire net957_c1;
wire net957;
wire net958_c1;
wire net958;
wire net959_c1;
wire net959;
wire net960_c1;
wire net960;
wire net961_c1;
wire net961;
wire net962_c1;
wire net962;
wire net963_c1;
wire net963;
wire net964_c1;
wire net964;
wire net965_c1;
wire net965;
wire net966_c1;
wire net966;
wire net967_c1;
wire net967;
wire net968_c1;
wire net968;
wire net969_c1;
wire net969;
wire net970_c1;
wire net970;
wire net971_c1;
wire net971;
wire net972_c1;
wire net972;
wire net973_c1;
wire net973;
wire net974_c1;
wire net974;
wire net975_c1;
wire net975;
wire net976_c1;
wire net976;
wire net977_c1;
wire net977;
wire net978_c1;
wire net978;
wire net979_c1;
wire net979;
wire net980_c1;
wire net980;
wire net981_c1;
wire net981;
wire net982_c1;
wire net982;
wire net983_c1;
wire net983;
wire net984_c1;
wire net984;
wire net985_c1;
wire net985;
wire net986_c1;
wire net986;
wire net987_c1;
wire net987;
wire net988_c1;
wire net988;
wire net989_c1;
wire net989;
wire net990_c1;
wire net990;
wire net991_c1;
wire net991;
wire net992_c1;
wire net992;
wire net993_c1;
wire net993;
wire net994_c1;
wire net994;
wire net995_c1;
wire net995;
wire net996_c1;
wire net996;
wire net997_c1;
wire net997;
wire net998_c1;
wire net998;
wire net999_c1;
wire net999;
wire net1000_c1;
wire net1000;
wire net1001_c1;
wire net1001;
wire net1002_c1;
wire net1002;
wire net1003_c1;
wire net1003;
wire net1004_c1;
wire net1004;
wire net1005_c1;
wire net1005;
wire net1006_c1;
wire net1006;
wire net1007_c1;
wire net1007;
wire net1008_c1;
wire net1008;
wire net1009_c1;
wire net1009;
wire net1010_c1;
wire net1010;
wire net1011_c1;
wire net1011;
wire net1012_c1;
wire net1012;
wire net1013_c1;
wire net1013;
wire net1014_c1;
wire net1014;
wire net1015_c1;
wire net1015;
wire net1016_c1;
wire net1016;
wire net1017_c1;
wire net1017;
wire net1018_c1;
wire net1018;
wire net1019_c1;
wire net1019;
wire net1020_c1;
wire net1020;
wire net1021_c1;
wire net1021;
wire net1022_c1;
wire net1022;
wire net1023_c1;
wire net1023;
wire net1024_c1;
wire net1024;
wire net1025_c1;
wire net1025;
wire net1026_c1;
wire net1026;
wire net1027_c1;
wire net1027;
wire net1028_c1;
wire net1028;
wire net1029_c1;
wire net1029;
wire net1030_c1;
wire net1030;
wire net1031_c1;
wire net1031;
wire net1032_c1;
wire net1032;
wire net1033_c1;
wire net1033;
wire net1034_c1;
wire net1034;
wire net1035_c1;
wire net1035;
wire net1036_c1;
wire net1036;
wire net1037_c1;
wire net1037;
wire net1038_c1;
wire net1038;
wire net1039_c1;
wire net1039;
wire net1040_c1;
wire net1040;
wire net1041_c1;
wire net1041;
wire net1042_c1;
wire net1042;
wire net1043_c1;
wire net1043;
wire net1044_c1;
wire net1044;
wire net1045_c1;
wire net1045;
wire net1046_c1;
wire net1046;
wire net1047_c1;
wire net1047;
wire net1048_c1;
wire net1048;
wire net1049_c1;
wire net1049;
wire net1050_c1;
wire net1050;
wire net1051_c1;
wire net1051;
wire net1052_c1;
wire net1052;
wire net1053_c1;
wire net1053;
wire net1054_c1;
wire net1054;
wire net1055_c1;
wire net1055;
wire net1056_c1;
wire net1056;
wire net1057_c1;
wire net1057;
wire net1058_c1;
wire net1058;
wire net1059_c1;
wire net1059;
wire net1060_c1;
wire net1060;
wire net1061_c1;
wire net1061;
wire net1062_c1;
wire net1062;
wire net1063_c1;
wire net1063;
wire net1064_c1;
wire net1064;
wire net1065_c1;
wire net1065;
wire net1066_c1;
wire net1066;
wire net1067_c1;
wire net1067;
wire net1068_c1;
wire net1068;
wire net1069_c1;
wire net1069;
wire net1070_c1;
wire net1070;
wire net1071_c1;
wire net1071;
wire net1072_c1;
wire net1072;
wire net1073_c1;
wire net1073;
wire net1074_c1;
wire net1074;
wire net1075_c1;
wire net1075;
wire net1076_c1;
wire net1076;
wire net1077_c1;
wire net1077;
wire net1078_c1;
wire net1078;
wire net1079_c1;
wire net1079;
wire net1080_c1;
wire net1080;
wire net1081_c1;
wire net1081;
wire net1082_c1;
wire net1082;
wire net1083_c1;
wire net1083;
wire net1084_c1;
wire net1084;
wire net1085_c1;
wire net1085;
wire net1086_c1;
wire net1086;
wire net1087_c1;
wire net1087;
wire net1088_c1;
wire net1088;
wire net1089_c1;
wire net1089;
wire net1090_c1;
wire net1090;
wire net1091_c1;
wire net1091;
wire net1092_c1;
wire net1092;
wire net1093_c1;
wire net1093;
wire net1094_c1;
wire net1094;
wire net1095_c1;
wire net1095;
wire net1096_c1;
wire net1096;
wire net1097_c1;
wire net1097;
wire net1098_c1;
wire net1098;
wire net1099_c1;
wire net1099;
wire net1100_c1;
wire net1100;
wire net1101_c1;
wire net1101;
wire net1102_c1;
wire net1102;
wire net1103_c1;
wire net1103;
wire net1104_c1;
wire net1104;
wire net1105_c1;
wire net1105;
wire net1106_c1;
wire net1106;
wire net1107_c1;
wire net1107;
wire net1108_c1;
wire net1108;
wire net1109_c1;
wire net1109;
wire net1110_c1;
wire net1110;
wire net1111_c1;
wire net1111;
wire net1112_c1;
wire net1112;
wire net1113_c1;
wire net1113;
wire net1114_c1;
wire net1114;
wire net1115_c1;
wire net1115;
wire net1116_c1;
wire net1116;
wire net1117_c1;
wire net1117;
wire net1118_c1;
wire net1118;
wire net1119_c1;
wire net1119;
wire net1120_c1;
wire net1120;
wire net1121_c1;
wire net1121;
wire net1122_c1;
wire net1122;
wire net1123_c1;
wire net1123;
wire net1124_c1;
wire net1124;
wire net1125_c1;
wire net1125;
wire net1126_c1;
wire net1126;
wire net1127_c1;
wire net1127;
wire net1128_c1;
wire net1128;
wire net1129_c1;
wire net1129;
wire net1130_c1;
wire net1130;
wire net1131_c1;
wire net1131;
wire net1132_c1;
wire net1132;
wire net1133_c1;
wire net1133;
wire net1134_c1;
wire net1134;
wire net1135_c1;
wire net1135;
wire net1136_c1;
wire net1136;
wire net1137_c1;
wire net1137;
wire net1138_c1;
wire net1138;
wire net1139_c1;
wire net1139;
wire net1140_c1;
wire net1140;
wire net1141_c1;
wire net1141;
wire net1142_c1;
wire net1142;
wire net1143_c1;
wire net1143;
wire net1144_c1;
wire net1144;
wire net1145_c1;
wire net1145;
wire net1146_c1;
wire net1146;
wire net1147_c1;
wire net1147;
wire net1148_c1;
wire net1148;
wire net1149_c1;
wire net1149;
wire net1150_c1;
wire net1150;
wire net1151_c1;
wire net1151;
wire net1152_c1;
wire net1152;
wire net1153_c1;
wire net1153;
wire net1154_c1;
wire net1154;
wire net1155_c1;
wire net1155;
wire net1156_c1;
wire net1156;
wire net1157_c1;
wire net1157;
wire net1158_c1;
wire net1158;
wire net1159_c1;
wire net1159;
wire net1160_c1;
wire net1160;
wire net1161_c1;
wire net1161;
wire net1162_c1;
wire net1162;
wire net1163_c1;
wire net1163;
wire net1164_c1;
wire net1164;
wire net1165_c1;
wire net1165;
wire net1166_c1;
wire net1166;
wire net1167_c1;
wire net1167;
wire net1168_c1;
wire net1168;
wire net1169_c1;
wire net1169;
wire net1170_c1;
wire net1170;
wire net1171_c1;
wire net1171;
wire net1172_c1;
wire net1172;
wire net1173_c1;
wire net1173;
wire net1174_c1;
wire net1174;
wire net1175_c1;
wire net1175;
wire net1176_c1;
wire net1176;
wire net1177_c1;
wire net1177;
wire net1178_c1;
wire net1178;
wire net1179_c1;
wire net1179;
wire net1180_c1;
wire net1180;
wire net1181_c1;
wire net1181;
wire net1182_c1;
wire net1182;
wire net1183_c1;
wire net1183;
wire net1184_c1;
wire net1184;
wire net1185_c1;
wire net1185;
wire net1186_c1;
wire net1186;
wire net1187_c1;
wire net1187;
wire net1188_c1;
wire net1188;
wire net1189_c1;
wire net1189;
wire net1190_c1;
wire net1190;
wire net1191_c1;
wire net1191;
wire net1192_c1;
wire net1192;
wire net1193_c1;
wire net1193;
wire net1194_c1;
wire net1194;
wire net1195_c1;
wire net1195;
wire net1196_c1;
wire net1196;
wire net1197_c1;
wire net1197;
wire net1198_c1;
wire net1198;
wire net1199_c1;
wire net1199;
wire net1200_c1;
wire net1200;
wire net1201_c1;
wire net1201;
wire net1202_c1;
wire net1202;
wire net1203_c1;
wire net1203;
wire net1204_c1;
wire net1204;
wire net1205_c1;
wire net1205;
wire net1206_c1;
wire net1206;
wire net1207_c1;
wire net1207;
wire net1208_c1;
wire net1208;
wire net1209_c1;
wire net1209;
wire net1210_c1;
wire net1210;
wire net1211_c1;
wire net1211;
wire net1212_c1;
wire net1212;
wire net1213_c1;
wire net1213;
wire net1214_c1;
wire net1214;
wire net1215_c1;
wire net1215;
wire net1216_c1;
wire net1216;
wire net1217_c1;
wire net1217;
wire net1218_c1;
wire net1218;
wire net1219_c1;
wire net1219;
wire net1220_c1;
wire net1220;
wire net1221_c1;
wire net1221;
wire net1222_c1;
wire net1222;
wire net1223_c1;
wire net1223;
wire net1224_c1;
wire net1224;
wire net1225_c1;
wire net1225;
wire net1226_c1;
wire net1226;
wire net1227_c1;
wire net1227;
wire net1228_c1;
wire net1228;
wire net1229_c1;
wire net1229;
wire net1230_c1;
wire net1230;
wire net1231_c1;
wire net1231;
wire net1232_c1;
wire net1232;
wire net1233_c1;
wire net1233;
wire net1234_c1;
wire net1234;
wire net1235_c1;
wire net1235;
wire net1236_c1;
wire net1236;
wire net1237_c1;
wire net1237;
wire net1238_c1;
wire net1238;
wire net1239_c1;
wire net1239;
wire net1240_c1;
wire net1240;
wire net1241_c1;
wire net1241;
wire net1242_c1;
wire net1242;
wire net1243_c1;
wire net1243;
wire net1244_c1;
wire net1244;
wire net1245_c1;
wire net1245;
wire net1246_c1;
wire net1246;
wire net1247_c1;
wire net1247;
wire net1248_c1;
wire net1248;
wire net1249_c1;
wire net1249;
wire net1250_c1;
wire net1250;
wire net1251_c1;
wire net1251;
wire net1252_c1;
wire net1252;
wire net1253_c1;
wire net1253;
wire net1254_c1;
wire net1254;
wire net1255_c1;
wire net1255;
wire net1256_c1;
wire net1256;
wire net1257_c1;
wire net1257;
wire net1258_c1;
wire net1258;
wire net1259_c1;
wire net1259;
wire net1260_c1;
wire net1260;
wire net1261_c1;
wire net1261;
wire net1262_c1;
wire net1262;
wire net1263_c1;
wire net1263;
wire net1264_c1;
wire net1264;
wire net1265_c1;
wire net1265;
wire net1266_c1;
wire net1266;
wire net1267_c1;
wire net1267;
wire net1268_c1;
wire net1268;
wire net1269_c1;
wire net1269;
wire net1270_c1;
wire net1270;
wire net1271_c1;
wire net1271;
wire net1272_c1;
wire net1272;
wire net1273_c1;
wire net1273;
wire net1274_c1;
wire net1274;
wire net1275_c1;
wire net1275;
wire net1276_c1;
wire net1276;
wire net1277_c1;
wire net1277;
wire net1278_c1;
wire net1278;
wire net1279_c1;
wire net1279;
wire net1280_c1;
wire net1280;
wire net1281_c1;
wire net1281;
wire net1282_c1;
wire net1282;
wire net1283_c1;
wire net1283;
wire net1284_c1;
wire net1284;
wire net1285_c1;
wire net1285;
wire net1286_c1;
wire net1286;
wire net1287_c1;
wire net1287;
wire net1288_c1;
wire net1288;
wire net1289_c1;
wire net1289;
wire net1290_c1;
wire net1290;
wire net1291_c1;
wire net1291;
wire net1292_c1;
wire net1292;
wire net1293_c1;
wire net1293;
wire net1294_c1;
wire net1294;
wire net1295_c1;
wire net1295;
wire net1296_c1;
wire net1296;
wire net1297_c1;
wire net1297;
wire net1298_c1;
wire net1298;
wire net1299_c1;
wire net1299;
wire net1300_c1;
wire net1300;
wire net1301_c1;
wire net1301;
wire net1302_c1;
wire net1302;
wire net1303_c1;
wire net1303;
wire net1304_c1;
wire net1304;
wire net1305_c1;
wire net1305;
wire net1306_c1;
wire net1306;
wire net1307_c1;
wire net1307;
wire net1308_c1;
wire net1308;
wire net1309_c1;
wire net1309;
wire net1310_c1;
wire net1310;
wire net1311_c1;
wire net1311;
wire net1312_c1;
wire net1312;
wire net1313_c1;
wire net1313;
wire net1314_c1;
wire net1314;
wire net1315_c1;
wire net1315;
wire net1316_c1;
wire net1316;
wire net1317_c1;
wire net1317;
wire net1318_c1;
wire net1318;
wire net1319_c1;
wire net1319;
wire net1320_c1;
wire net1320;
wire net1321_c1;
wire net1321;
wire net1322_c1;
wire net1322;
wire net1323_c1;
wire net1323;
wire net1324_c1;
wire net1324;
wire net1325_c1;
wire net1325;
wire net1326_c1;
wire net1326;
wire net1327_c1;
wire net1327;
wire net1328_c1;
wire net1328;
wire net1329_c1;
wire net1329;
wire net1330_c1;
wire net1330;
wire net1331_c1;
wire net1331;
wire net1332_c1;
wire net1332;
wire net1333_c1;
wire net1333;
wire net1334_c1;
wire net1334;
wire net1335_c1;
wire net1335;
wire net1336_c1;
wire net1336;
wire net1337_c1;
wire net1337;
wire net1338_c1;
wire net1338;
wire net1339_c1;
wire net1339;
wire net1340_c1;
wire net1340;
wire net1341_c1;
wire net1341;
wire net1342_c1;
wire net1342;
wire net1343_c1;
wire net1343;
wire net1344_c1;
wire net1344;
wire net1345_c1;
wire net1345;
wire net1346_c1;
wire net1346;
wire net1347_c1;
wire net1347;
wire net1348_c1;
wire net1348;
wire net1349_c1;
wire net1349;
wire net1350_c1;
wire net1350;
wire net1351_c1;
wire net1351;
wire net1352_c1;
wire net1352;
wire net1353_c1;
wire net1353;
wire net1354_c1;
wire net1354;
wire net1355_c1;
wire net1355;
wire net1356_c1;
wire net1356;
wire net1357_c1;
wire net1357;
wire net1358_c1;
wire net1358;
wire net1359_c1;
wire net1359;
wire GCLK_Pad;
wire net1360;
wire net1361_c1;
wire net1361;
wire net1362_c1;
wire net1362;
wire net1363_c1;
wire net1363;

DFFT DFFT_295__FPB_n751(net1266,net467,net477_c1);
DFFT DFFT_287__FPB_n743(net765,net468,net478_c1);
DFFT DFFT_279__FPB_n735(net764,net1362,net479_c1);
DFFT DFFT_199__FPB_n655(net763,net471,net485_c1);
DFFT DFFT_296__FPB_n752(net762,net477,net488_c1);
DFFT DFFT_288__FPB_n744(net761,net478,net489_c1);
DFFT DFFT_297__FPB_n753(net1060,net488,net498_c1);
DFFT DFFT_289__FPB_n745(net1042,net489,net499_c1);
DFFT DFFT_306_state_obs3(net1267,net497,net550_c1);
DFFT DFFT_298__FPB_n754(net760,net498,net507_c1);
XOR2T XOR2T_36_n60(net759,net337,net388,net11_c1);
XOR2T XOR2T_45_n69(net758,net285,net1363,net56_c1);
XOR2T XOR2T_55_n79(net757,net173,net495,net62_c1);
AND2T AND2T_101_n125(net756,net378,net544,net96_c1);
AND2T AND2T_110_n134(net755,net153,net194,net101_c1);
AND2T AND2T_103_n127(net754,net102,net276,net107_c1);
AND2T AND2T_104_n128(net753,net202,net546,net113_c1);
AND2T AND2T_121_n145(net1322,net105,net426,net116_c1);
AND2T AND2T_113_n137(net752,net358,net179,net117_c1);
AND2T AND2T_105_n129(net751,net252,net417,net118_c1);
AND2T AND2T_106_n130(net1100,net364,net418,net81_c1);
AND2T AND2T_122_n146(net750,net151,net438,net121_c1);
AND2T AND2T_114_n138(net749,net17,net28,net122_c1);
AND2T AND2T_123_n147(net748,net390,net453,net125_c1);
AND2T AND2T_132_n156(net747,net229,net425,net128_c1);
AND2T AND2T_124_n148(net1210,net132,net462,net129_c1);
AND2T AND2T_140_n176(net746,net361,net352,net138_c1);
AND2T AND2T_109_n133(net745,net226,net424,net95_c1);
AND2T AND2T_133_n157(net744,net335,net437,net131_c1);
AND2T AND2T_141_n177(net743,net319,net452,net139_c1);
AND2T AND2T_143_n179(net1024,net13,net311,net141_c1);
AND2T AND2T_128_n152(net742,net239,net484,net110_c1);
AND2T AND2T_144_n180(net741,net3,net461,net127_c1);
AND2T AND2T_129_n153(net740,net110,net104,net115_c1);
AND2T AND2T_145_n181(net1025,net185,net472,net130_c1);
AND2T AND2T_146_n182(net739,net374,net367,net133_c1);
AND2T AND2T_139_n163(net738,net114,net445,net123_c1);
AND2T AND2T_9_n33(net737,net354,net421,net4_c1);
NOTT NOTT_8_n32(net736,net336,net2_c1);
AND2T AND2T_10_n34(net735,net231,net429,net7_c1);
AND2T AND2T_11_n35(net1340,net363,net441,net10_c1);
AND2T AND2T_12_n36(net1276,net240,net457,net14_c1);
AND2T AND2T_21_n45(net734,net323,net341,net17_c1);
AND2T AND2T_13_n37(net733,net375,net389,net18_c1);
AND2T AND2T_22_n46(net732,net324,net342,net22_c1);
AND2T AND2T_15_n39(net731,net313,net466,net28_c1);
AND2T AND2T_16_n40(net1136,net296,net476,net1_c1);
AND2T AND2T_32_n56(net730,net170,net448,net32_c1);
AND2T AND2T_24_n48(net1232,net181,net486,net33_c1);
AND2T AND2T_33_n57(net729,net212,net175,net37_c1);
AND2T AND2T_25_n49(net728,net204,net428,net38_c1);
AND2T AND2T_26_n50(net904,net334,net292,net5_c1);
AND2T AND2T_18_n42(net727,net188,net303,net6_c1);
AND2T AND2T_27_n51(net1248,net222,net434,net8_c1);
AND2T AND2T_51_n75(net726,net298,net447,net46_c1);
AND2T AND2T_43_n67(net840,net31,net475,net47_c1);
AND2T AND2T_35_n59(net725,net187,net456,net48_c1);
AND2T AND2T_28_n52(net724,net230,net267,net12_c1);
AND2T AND2T_52_n76(net788,net343,net455,net51_c1);
AND2T AND2T_44_n68(net1016,net56,net496,net52_c1);
AND2T AND2T_29_n53(net723,net307,net440,net16_c1);
AND2T AND2T_61_n85(net722,net210,net284,net54_c1);
AND2T AND2T_53_n77(net721,net51,net464,net55_c1);
AND2T AND2T_46_n70(net720,net366,net24,net19_c1);
AND2T AND2T_54_n78(net719,net221,net485,net59_c1);
AND2T AND2T_39_n63(net912,net297,net203,net25_c1);
AND2T AND2T_71_n95(net718,net370,net174,net60_c1);
AND2T AND2T_63_n87(net717,net58,net494,net61_c1);
AND2T AND2T_56_n80(net1084,net272,net505,net29_c1);
AND2T AND2T_48_n72(net716,net35,net439,net30_c1);
AND2T AND2T_72_n96(net715,net277,net520,net63_c1);
AND2T AND2T_64_n88(net714,net161,net504,net64_c1);
AND2T AND2T_57_n81(net713,net247,net514,net34_c1);
AND2T AND2T_73_n97(net804,net263,net526,net65_c1);
AND2T AND2T_66_n90(net712,net196,net355,net39_c1);
AND2T AND2T_67_n91(net711,net348,net227,net44_c1);
AND2T AND2T_68_n92(net710,net44,net305,net49_c1);
DFFT DFFT_292_state_obs1(net986,net515,net548_c1);
OR2T OR2T_30_n54(net876,net381,net349,net21_c1);
OR2T OR2T_31_n55(net709,net21,net27,net26_c1);
OR2T OR2T_23_n47(net877,net369,net327,net27_c1);
OR2T OR2T_42_n66(net708,net359,net317,net42_c1);
OR2T OR2T_34_n58(net707,net344,net386,net43_c1);
OR2T OR2T_60_n84(net706,net45,net454,net50_c1);
OR2T OR2T_37_n61(net805,net43,net465,net15_c1);
OR2T OR2T_38_n62(net705,net15,net26,net20_c1);
OR2T OR2T_70_n94(net704,net53,net66,net57_c1);
OR2T OR2T_62_n86(net703,net228,net463,net58_c1);
OR2T OR2T_65_n89(net702,net273,net259,net66_c1);
OR2T OR2T_58_n82(net701,net302,net521,net40_c1);
OR2T OR2T_74_n98(net700,net65,net63,net67_c1);
OR2T OR2T_59_n83(net699,net34,net29,net45_c1);
OR2T OR2T_75_n99(net698,net67,net57,net68_c1);
OR2T OR2T_69_n93(net905,net49,net275,net53_c1);
DFFT DFFT_285_state_obs0(net697,net449,net547_c1);
NOTT NOTT_20_n44(net696,net254,net13_c1);
NOTT NOTT_14_n38(net695,net353,net23_c1);
NOTT NOTT_40_n64(net694,net350,net31_c1);
NOTT NOTT_17_n41(net693,net392,net3_c1);
NOTT NOTT_41_n65(net692,net331,net36_c1);
NOTT NOTT_50_n74(net691,net356,net41_c1);
NOTT NOTT_19_n43(net690,net264,net9_c1);
NOTT NOTT_47_n71(net689,net52,net24_c1);
NOTT NOTT_49_n73(net688,net20,net35_c1);
OR2T OR2T_100_n124(net1233,net209,net9,net91_c1);
OR2T OR2T_102_n126(net687,net278,net219,net102_c1);
OR2T OR2T_111_n135(net913,net101,net148,net106_c1);
OR2T OR2T_112_n136(net686,net106,net427,net112_c1);
OR2T OR2T_130_n154(net1118,net150,net154,net120_c1);
OR2T OR2T_107_n131(net1156,net81,net113,net85_c1);
OR2T OR2T_131_n155(net1137,net120,net115,net124_c1);
OR2T OR2T_115_n139(net1192,net287,net283,net126_c1);
OR2T OR2T_116_n140(net1193,net126,net165,net89_c1);
OR2T OR2T_108_n132(net685,net85,net420,net90_c1);
OR2T OR2T_117_n141(net684,net89,net112,net94_c1);
OR2T OR2T_125_n149(net683,net164,net159,net132_c1);
OR2T OR2T_126_n150(net1211,net129,net473,net99_c1);
OR2T OR2T_118_n142(net682,net94,net90,net100_c1);
OR2T OR2T_134_n158(net1128,net131,net128,net134_c1);
OR2T OR2T_127_n151(net681,net281,net376,net104_c1);
OR2T OR2T_119_n143(net680,net387,net433,net105_c1);
OR2T OR2T_135_n159(net679,net134,net124,net136_c1);
OR2T OR2T_136_n160(net678,net136,net99,net109_c1);
OR2T OR2T_137_n161(net677,net261,net446,net114_c1);
DFFT DFFT_299_state_obs2(net676,net507,net549_c1);
AND2T AND2T_80_n104(net675,net72,net531,net77_c1);
AND2T AND2T_81_n105(net674,net84,net513,net80_c1);
AND2T AND2T_90_n114(net822,net330,net365,net83_c1);
AND2T AND2T_91_n115(net673,net146,net530,net87_c1);
AND2T AND2T_83_n107(net672,net225,net93,net88_c1);
AND2T AND2T_92_n116(net671,net220,net540,net92_c1);
AND2T AND2T_84_n108(net670,net262,net379,net93_c1);
AND2T AND2T_85_n109(net669,net309,net314,net98_c1);
AND2T AND2T_86_n110(net1119,net98,net245,net71_c1);
AND2T AND2T_87_n111(net668,net271,net320,net73_c1);
AND2T AND2T_98_n122(net1006,net75,net539,net82_c1);
AND2T AND2T_99_n123(net667,net91,net541,net86_c1);
DFFT DFFT_200__FPB_n656(net666,net253,net495_c1);
DFFT DFFT_201__FPB_n657(net665,net62,net505_c1);
DFFT DFFT_155__PIPL_n209(net664,net4,net399_c1);
DFFT DFFT_210__FPB_n666(net663,net195,net512_c1);
DFFT DFFT_202__FPB_n658(net662,net40,net514_c1);
DFFT DFFT_211__FPB_n667(net1085,net512,net520_c1);
DFFT DFFT_203__FPB_n659(net661,net351,net521_c1);
DFFT DFFT_156__PIPL_n210(net660,net7,net396_c1);
DFFT DFFT_204__FPB_n660(net659,net55,net454_c1);
DFFT DFFT_300__FPB_n756(net1358,net398,net522_c1);
DFFT DFFT_220__FPB_n676(net950,net519,net524_c1);
DFFT DFFT_212__FPB_n668(net658,net393,net526_c1);
DFFT DFFT_205__FPB_n661(net841,net54,net463_c1);
DFFT DFFT_301__FPB_n757(net1359,net522,net527_c1);
DFFT DFFT_221__FPB_n677(net978,net524,net531_c1);
DFFT DFFT_213__FPB_n669(net657,net61,net532_c1);
DFFT DFFT_157__PIPL_n211(net1341,net10,net397_c1);
DFFT DFFT_214__FPB_n670(net656,net50,net474_c1);
DFFT DFFT_206__FPB_n662(net655,net180,net470_c1);
DFFT DFFT_302__FPB_n758(net1284,net527,net533_c1);
DFFT DFFT_230__FPB_n686(net654,net322,net535_c1);
DFFT DFFT_222__FPB_n678(net653,net238,net536_c1);
DFFT DFFT_215__FPB_n671(net652,net74,net481_c1);
DFFT DFFT_207__FPB_n663(net651,net470,net482_c1);
DFFT DFFT_303__FPB_n759(net1285,net533,net537_c1);
DFFT DFFT_231__FPB_n687(net650,net535,net540_c1);
DFFT DFFT_223__FPB_n679(net823,net536,net538_c1);
DFFT DFFT_160__FBL_n616(net1007,net299,net405_c1);
OR2T OR2T_76_n100(net649,net68,net532,net69_c1);
DFFT DFFT_158__PIPL_n212(net648,net14,net398_c1);
OR2T OR2T_77_n101(net789,net69,net474,net70_c1);
OR2T OR2T_93_n117(net647,net290,net87,net97_c1);
OR2T OR2T_78_n102(net646,net70,net382,net72_c1);
DFFT DFFT_152__FPB_n206(net645,net326,net414_c1);
OR2T OR2T_94_n118(net644,net97,net79,net103_c1);
DFFT DFFT_304__FPB_n760(net643,net537,net487_c1);
DFFT DFFT_224__FPB_n680(net642,net538,net492_c1);
DFFT DFFT_216__FPB_n672(net641,net481,net493_c1);
DFFT DFFT_208__FPB_n664(net640,net482,net494_c1);
OR2T OR2T_95_n119(net639,net80,net542,net108_c1);
DFFT DFFT_240__FPB_n696(net1017,net249,net541_c1);
DFFT DFFT_232__FPB_n688(net638,net103,net542_c1);
OR2T OR2T_96_n120(net637,net108,net258,net75_c1);
OR2T OR2T_88_n112(net894,net73,net71,net76_c1);
OR2T OR2T_89_n113(net636,net76,net525,net79_c1);
DFFT DFFT_161__FBL_n617(net1314,net300,net407_c1);
DFFT DFFT_153__FPB_n207(net1157,net201,net415_c1);
DFFT DFFT_305__FPB_n761(net635,net487,net497_c1);
DFFT DFFT_225__FPB_n681(net634,net492,net502_c1);
DFFT DFFT_217__FPB_n673(net633,net493,net503_c1);
DFFT DFFT_209__FPB_n665(net632,net377,net504_c1);
DFFT DFFT_241__FPB_n697(net860,net372,net544_c1);
DFFT DFFT_233__FPB_n689(net631,net78,net543_c1);
DFFT DFFT_170__FBL_n626(net630,net310,net409_c1);
DFFT DFFT_162__FBL_n618(net629,net279,net410_c1);
DFFT DFFT_154__FPB_n208(net628,net207,net416_c1);
DFFT DFFT_250__FPB_n706(net627,net111,net436_c1);
DFFT DFFT_234__FPB_n690(net1052,net543,net510_c1);
DFFT DFFT_226__FPB_n682(net626,net502,net513_c1);
DFFT DFFT_218__FPB_n674(net625,net503,net511_c1);
DFFT DFFT_242__FPB_n698(net624,net200,net545_c1);
DFFT DFFT_171__FBL_n627(net1249,net147,net411_c1);
DFFT DFFT_163__FBL_n619(net623,net158,net412_c1);
DFFT DFFT_251__FPB_n707(net622,net436,net443_c1);
DFFT DFFT_235__FPB_n691(net1053,net510,net517_c1);
DFFT DFFT_227__FPB_n683(net832,net88,net518_c1);
DFFT DFFT_219__FPB_n675(net621,net511,net519_c1);
DFFT DFFT_243__FPB_n699(net1166,net545,net546_c1);
DFFT DFFT_164__FBL_n620(net620,net172,net400_c1);
DFFT DFFT_172__FBL_n628(net1323,net178,net413_c1);
DFFT DFFT_244__FPB_n700(net619,net383,net417_c1);
DFFT DFFT_260__FPB_n716(net618,net442,net453_c1);
DFFT DFFT_252__FPB_n708(net617,net443,net451_c1);
DFFT DFFT_180__FPB_n636(net616,net444,net457_c1);
DFFT DFFT_236__FPB_n692(net615,net517,net523_c1);
DFFT DFFT_228__FPB_n684(net833,net518,net525_c1);
DFFT DFFT_165__FBL_n621(net614,net171,net401_c1);
DFFT DFFT_245__FPB_n701(net1101,net157,net418_c1);
DFFT DFFT_261__FPB_n717(net1202,net125,net462_c1);
DFFT DFFT_253__FPB_n709(net1350,net451,net459_c1);
DFFT DFFT_181__FPB_n637(net613,net270,net466_c1);
DFFT DFFT_173__FPB_n629(net612,net391,net460_c1);
DFFT DFFT_237__FPB_n693(net611,net523,net529_c1);
DFFT DFFT_229__FPB_n685(net610,net83,net530_c1);
DFFT DFFT_166__FBL_n622(net609,net152,net402_c1);
DFFT DFFT_254__FPB_n710(net1351,net459,net419_c1);
DFFT DFFT_246__FPB_n702(net608,net107,net420_c1);
DFFT DFFT_174__FPB_n630(net979,net460,net421_c1);
DFFT DFFT_270__FPB_n726(net607,net458,net469_c1);
DFFT DFFT_262__FPB_n718(net1203,net121,net473_c1);
DFFT DFFT_190__FPB_n646(net895,net42,net475_c1);
DFFT DFFT_182__FPB_n638(net606,net160,net476_c1);
DFFT DFFT_238__FPB_n694(net605,net529,net534_c1);
DFFT DFFT_167__FBL_n623(net951,net280,net403_c1);
DFFT DFFT_159__FBL_n615(net604,net286,net404_c1);
SPLITT Split_310_n766(net149,net207_c1,net338_c1);
SPLITT Split_311_n767(net2,net215_c1,net347_c1);
SPLITT Split_312_n768(net347,net231_c1,net354_c1);
SPLITT Split_320_n776(net206,net226_c1,net355_c1);
SPLITT Split_400_n856(net339,net227_c1,net356_c1);
SPLITT Split_313_n769(net215,net240_c1,net363_c1);
SPLITT Split_321_n777(net22,net237_c1,net364_c1);
SPLITT Split_401_n857(net214,net238_c1,net365_c1);
SPLITT Split_314_n770(net23,net177_c1,net306_c1);
SPLITT Split_322_n778(net237,net247_c1,net369_c1);
SPLITT Split_330_n786(net236,net245_c1,net370_c1);
SPLITT Split_402_n858(net415,net242_c1,net371_c1);
SPLITT Split_410_n866(net405,net243_c1,net372_c1);
SPLITT Split_307_n763(net0,net183_c1,net312_c1);
SPLITT Split_315_n771(net306,net188_c1,net313_c1);
SPLITT Split_323_n779(net33,net251_c1,net376_c1);
SPLITT Split_331_n787(net12,net249_c1,net377_c1);
SPLITT Split_403_n859(net371,net252_c1,net378_c1);
SPLITT Split_411_n867(net243,net253_c1,net379_c1);
SPLITT Split_308_n764(net312,net192_c1,net318_c1);
SPLITT Split_316_n772(net177,net193_c1,net319_c1);
SPLITT Split_324_n780(net251,net194_c1,net320_c1);
SPLITT Split_404_n860(net242,net191_c1,net321_c1);
SPLITT Split_332_n788(net16,net259_c1,net381_c1);
SPLITT Split_340_n796(net373,net258_c1,net382_c1);
SPLITT Split_412_n868(net407,net256_c1,net383_c1);
SPLITT Split_420_n876(net403,net255_c1,net384_c1);
SPLITT Split_309_n765(net183,net201_c1,net326_c1);
SPLITT Split_317_n773(net1,net202_c1,net327_c1);
SPLITT Split_325_n781(net38,net199_c1,net328_c1);
SPLITT Split_405_n861(net416,net197_c1,net329_c1);
SPLITT Split_333_n789(net32,net263_c1,net386_c1);
SPLITT Split_341_n797(net248,net261_c1,net387_c1);
SPLITT Split_413_n869(net256,net262_c1,net388_c1);
SPLITT Split_421_n877(net384,net264_c1,net389_c1);
SPLITT Split_350_n806(net156,net158_c1,net286_c1);
SPLITT Split_318_n774(net6,net206_c1,net333_c1);
SPLITT Split_326_n782(net328,net212_c1,net334_c1);
SPLITT Split_334_n790(net37,net208_c1,net335_c1);
SPLITT Split_406_n862(net329,net213_c1,net336_c1);
SPLITT Split_414_n870(net410,net211_c1,net337_c1);
SPLITT Split_342_n798(net41,net266_c1,net390_c1);
SPLITT Split_422_n878(net255,net265_c1,net391_c1);
SPLITT Split_430_n886(net385,net267_c1,net392_c1);
SPLITT Split_351_n807(net92,net165_c1,net290_c1);
SPLITT Split_319_n775(net333,net221_c1,net342_c1);
SPLITT Split_327_n783(net199,net219_c1,net343_c1);
SPLITT Split_335_n791(net208,net220_c1,net344_c1);
SPLITT Split_407_n863(net197,net218_c1,net345_c1);
SPLITT Split_415_n871(net412,net217_c1,net346_c1);
SPLITT Split_343_n799(net46,net269_c1,net393_c1);
SPLITT Split_423_n879(net409,net268_c1,net394_c1);
SPLITT Split_431_n887(net260,net270_c1,net395_c1);
SPLITT Split_344_n800(net269,net145_c1,net271_c1);
SPLITT Split_352_n808(net82,net169_c1,net294_c1);
SPLITT Split_360_n816(net116,net168_c1,net295_c1);
SPLITT Split_328_n784(net5,net229_c1,net349_c1);
SPLITT Split_336_n792(net25,net228_c1,net350_c1);
SPLITT Split_408_n864(net404,net223_c1,net351_c1);
SPLITT Split_416_n872(net217,net224_c1,net352_c1);
SPLITT Split_424_n880(net394,net230_c1,net353_c1);
SPLITT Split_345_n801(net59,net146_c1,net272_c1);
SPLITT Split_353_n809(net294,net172_c1,net299_c1);
SPLITT Split_361_n817(net295,net171_c1,net300_c1);
SPLITT Split_329_n785(net8,net236_c1,net358_c1);
SPLITT Split_337_n793(net36,net239_c1,net359_c1);
SPLITT Split_409_n865(net223,net233_c1,net360_c1);
SPLITT Split_417_n873(net400,net235_c1,net361_c1);
SPLITT Split_425_n881(net268,net234_c1,net362_c1);
DFFT DFFT_255__FPB_n711(net603,net419,net422_c1);
DFFT DFFT_247__FPB_n703(net602,net163,net424_c1);
DFFT DFFT_175__FPB_n631(net1061,net380,net423_c1);
SPLITT Split_346_n802(net64,net148_c1,net273_c1);
SPLITT Split_354_n810(net169,net147_c1,net274_c1);
DFFT DFFT_271__FPB_n727(net601,net469,net480_c1);
DFFT DFFT_263__FPB_n719(net600,net18,net484_c1);
DFFT DFFT_191__FPB_n647(net599,net193,net483_c1);
DFFT DFFT_183__FPB_n639(net598,net234,net486_c1);
SPLITT Split_362_n818(net168,net178_c1,net304_c1);
SPLITT Split_370_n826(net167,net179_c1,net305_c1);
DFFT DFFT_239__FPB_n695(net597,net534,net539_c1);
SPLITT Split_338_n794(net47,net246_c1,net366_c1);
SPLITT Split_418_n874(net401,net244_c1,net367_c1);
SPLITT Split_426_n882(net411,net241_c1,net368_c1);
SPLITT Split_347_n803(net39,net151_c1,net275_c1);
SPLITT Split_355_n811(net86,net150_c1,net276_c1);
SPLITT Split_363_n819(net123,net184_c1,net310_c1);
SPLITT Split_371_n827(net140,net185_c1,net311_c1);
SPLITT Split_339_n795(net30,net248_c1,net373_c1);
SPLITT Split_419_n875(net402,net250_c1,net374_c1);
SPLITT Split_427_n883(net368,net254_c1,net375_c1);
SPLITT Split_348_n804(net60,net154_c1,net277_c1);
SPLITT Split_356_n812(net96,net153_c1,net278_c1);
SPLITT Split_364_n820(net184,net152_c1,net279_c1);
SPLITT Split_372_n828(net141,net190_c1,net316_c1);
SPLITT Split_380_n836(net176,net196_c1,net317_c1);
SPLITT Split_428_n884(net241,net257_c1,net380_c1);
SPLITT Split_349_n805(net77,net156_c1,net280_c1);
SPLITT Split_357_n813(net118,net157_c1,net281_c1);
SPLITT Split_365_n821(net138,net155_c1,net282_c1);
SPLITT Split_373_n829(net316,net203_c1,net324_c1);
SPLITT Split_381_n837(net133,net198_c1,net325_c1);
SPLITT Split_429_n885(net413,net260_c1,net385_c1);
SPLITT Split_358_n814(net117,net159_c1,net283_c1);
SPLITT Split_366_n822(net282,net160_c1,net284_c1);
SPLITT Split_374_n830(net190,net161_c1,net285_c1);
SPLITT Split_382_n838(net325,net210_c1,net331_c1);
SPLITT Split_390_n846(net142,net205_c1,net332_c1);
SPLITT Split_359_n815(net122,net164_c1,net287_c1);
SPLITT Split_367_n823(net155,net163_c1,net288_c1);
SPLITT Split_375_n831(net127,net162_c1,net289_c1);
SPLITT Split_383_n839(net198,net216_c1,net340_c1);
SPLITT Split_391_n847(net332,net222_c1,net341_c1);
SPLITT Split_368_n824(net139,net167_c1,net291_c1);
SPLITT Split_376_n832(net289,net170_c1,net292_c1);
SPLITT Split_384_n840(net135,net166_c1,net293_c1);
SPLITT Split_392_n848(net205,net225_c1,net348_c1);
SPLITT Split_369_n825(net291,net175_c1,net296_c1);
SPLITT Split_377_n833(net162,net174_c1,net297_c1);
SPLITT Split_385_n841(net293,net173_c1,net298_c1);
SPLITT Split_393_n849(net143,net232_c1,net357_c1);
SPLITT Split_378_n834(net130,net176_c1,net301_c1);
SPLITT Split_386_n842(net166,net180_c1,net302_c1);
SPLITT Split_394_n850(net357,net181_c1,net303_c1);
SPLITT Split_379_n835(net301,net187_c1,net307_c1);
SPLITT Split_387_n843(net137,net182_c1,net308_c1);
SPLITT Split_395_n851(net232,net186_c1,net309_c1);
SPLITT Split_388_n844(net308,net195_c1,net314_c1);
SPLITT Split_396_n852(net144,net189_c1,net315_c1);
SPLITT Split_389_n845(net182,net200_c1,net322_c1);
SPLITT Split_397_n853(net315,net204_c1,net323_c1);
SPLITT Split_398_n854(net189,net209_c1,net330_c1);
SPLITT Split_399_n855(net414,net214_c1,net339_c1);
NOTT NOTT_120_n144(net1277,net218,net111_c1);
DFFT DFFT_168__FBL_n624(net596,net274,net406_c1);
NOTT NOTT_142_n178(net595,net224,net140_c1);
NOTT NOTT_150_n198(net1304,net1361,net143_c1);
NOTT NOTT_151_n199(net594,net406,net144_c1);
NOTT NOTT_138_n162(net593,net338,net119_c1);
NOTT NOTT_147_n183(net592,net318,net135_c1);
NOTT NOTT_148_n184(net591,net192,net137_c1);
NOTT NOTT_149_n197(net934,net346,net142_c1);
DFFT DFFT_264__FPB_n720(net1129,net266,net425_c1);
DFFT DFFT_256__FPB_n712(net590,net422,net426_c1);
DFFT DFFT_248__FPB_n704(net589,net95,net427_c1);
DFFT DFFT_184__FPB_n640(net935,net265,net428_c1);
DFFT DFFT_176__FPB_n632(net588,net423,net429_c1);
DFFT DFFT_280__FPB_n736(net587,net479,net490_c1);
DFFT DFFT_272__FPB_n728(net586,net480,net491_c1);
DFFT DFFT_192__FPB_n648(net585,net483,net496_c1);
DFFT DFFT_169__FBL_n625(net1305,net304,net408_c1);
DFFT DFFT_265__FPB_n721(net1167,net191,net430_c1);
DFFT DFFT_257__FPB_n713(net584,net321,net431_c1);
DFFT DFFT_249__FPB_n705(net1315,net100,net433_c1);
DFFT DFFT_185__FPB_n641(net583,net257,net434_c1);
DFFT DFFT_177__FPB_n633(net582,net395,net432_c1);
DFFT DFFT_281__FPB_n737(net581,net490,net500_c1);
DFFT DFFT_273__FPB_n729(net580,net491,net501_c1);
DFFT DFFT_193__FPB_n649(net579,net186,net506_c1);
DFFT DFFT_274__FPB_n730(net578,net501,net435_c1);
DFFT DFFT_266__FPB_n722(net1174,net430,net437_c1);
DFFT DFFT_258__FPB_n714(net1175,net431,net438_c1);
DFFT DFFT_194__FPB_n650(net577,net19,net439_c1);
DFFT DFFT_186__FPB_n642(net576,net340,net440_c1);
DFFT DFFT_178__FPB_n634(net575,net432,net441_c1);
DFFT DFFT_290__FPB_n746(net1043,net499,net508_c1);
DFFT DFFT_282__FPB_n738(net574,net500,net509_c1);
DFFT DFFT_275__FPB_n731(net573,net435,net445_c1);
DFFT DFFT_267__FPB_n723(net572,net109,net446_c1);
DFFT DFFT_259__FPB_n715(net571,net211,net442_c1);
DFFT DFFT_195__FPB_n651(net570,net360,net447_c1);
DFFT DFFT_187__FPB_n643(net569,net288,net448_c1);
DFFT DFFT_179__FPB_n635(net568,net362,net444_c1);
DFFT DFFT_291__FPB_n747(net987,net508,net515_c1);
DFFT DFFT_283__FPB_n739(net968,net509,net516_c1);
NOTT NOTT_82_n106(net567,net246,net84_c1);
DFFT DFFT_284__FPB_n740(net969,net516,net449_c1);
DFFT DFFT_276__FPB_n732(net566,net244,net452_c1);
DFFT DFFT_268__FPB_n724(net565,net119,net450_c1);
DFFT DFFT_196__FPB_n652(net564,net216,net455_c1);
DFFT DFFT_188__FPB_n644(net563,net11,net456_c1);
NOTT NOTT_79_n103(net562,net213,net74_c1);
NOTT NOTT_97_n121(net561,net345,net78_c1);
DFFT DFFT_277__FPB_n733(net560,net250,net461_c1);
DFFT DFFT_269__FPB_n725(net559,net450,net458_c1);
DFFT DFFT_197__FPB_n653(net558,net145,net464_c1);
DFFT DFFT_189__FPB_n645(net861,net48,net465_c1);
DFFT DFFT_293__FPB_n749(net557,net397,net528_c1);
DFFT DFFT_294__FPB_n750(net556,net528,net467_c1);
DFFT DFFT_286__FPB_n742(net555,net396,net468_c1);
DFFT DFFT_278__FPB_n734(net554,net235,net472_c1);
DFFT DFFT_198__FPB_n654(net553,net233,net471_c1);
SPLITT SplitCLK_4_300(net1357,net1358_c1,net1359_c1);
SPLITT SplitCLK_4_301(net1352,net1357_c1,net1356_c1);
SPLITT SplitCLK_6_302(net1353,net1354_c1,net1355_c1);
SPLITT SplitCLK_6_303(net1342,net1352_c1,net1353_c1);
SPLITT SplitCLK_4_304(net1349,net1350_c1,net1351_c1);
SPLITT SplitCLK_0_305(net1344,net1349_c1,net1348_c1);
SPLITT SplitCLK_2_306(net1345,net1347_c1,net1346_c1);
SPLITT SplitCLK_6_307(net1343,net1344_c1,net1345_c1);
SPLITT SplitCLK_4_308(net1324,net1343_c1,net1342_c1);
SPLITT SplitCLK_4_309(net1339,net1341_c1,net1340_c1);
SPLITT SplitCLK_4_310(net1334,net1339_c1,net1338_c1);
SPLITT SplitCLK_2_311(net1335,net1336_c1,net1337_c1);
SPLITT SplitCLK_6_312(net1326,net1334_c1,net1335_c1);
SPLITT SplitCLK_0_313(net1328,net1333_c1,net1332_c1);
SPLITT SplitCLK_2_314(net1329,net1330_c1,net1331_c1);
SPLITT SplitCLK_4_315(net1327,net1329_c1,net1328_c1);
SPLITT SplitCLK_2_316(net1325,net1327_c1,net1326_c1);
SPLITT SplitCLK_6_317(net1286,net1324_c1,net1325_c1);
SPLITT SplitCLK_4_318(net1321,net1322_c1,net1323_c1);
SPLITT SplitCLK_4_319(net1316,net1321_c1,net1320_c1);
SPLITT SplitCLK_2_320(net1317,net1318_c1,net1319_c1);
SPLITT SplitCLK_6_321(net1306,net1316_c1,net1317_c1);
SPLITT SplitCLK_4_322(net1313,net1314_c1,net1315_c1);
SPLITT SplitCLK_4_323(net1308,net1312_c1,net1313_c1);
SPLITT SplitCLK_2_324(net1309,net1310_c1,net1311_c1);
SPLITT SplitCLK_4_325(net1307,net1309_c1,net1308_c1);
SPLITT SplitCLK_4_326(net1288,net1306_c1,net1307_c1);
SPLITT SplitCLK_4_327(net1303,net1304_c1,net1305_c1);
SPLITT SplitCLK_4_328(net1298,net1303_c1,net1302_c1);
SPLITT SplitCLK_6_329(net1299,net1300_c1,net1301_c1);
SPLITT SplitCLK_6_330(net1290,net1298_c1,net1299_c1);
SPLITT SplitCLK_4_331(net1292,net1296_c1,net1297_c1);
SPLITT SplitCLK_6_332(net1293,net1295_c1,net1294_c1);
SPLITT SplitCLK_4_333(net1291,net1293_c1,net1292_c1);
SPLITT SplitCLK_2_334(net1289,net1291_c1,net1290_c1);
SPLITT SplitCLK_4_335(net1287,net1289_c1,net1288_c1);
SPLITT SplitCLK_0_336(net1212,net1286_c1,net1287_c1);
SPLITT SplitCLK_4_337(net1283,net1285_c1,net1284_c1);
SPLITT SplitCLK_4_338(net1278,net1283_c1,net1282_c1);
SPLITT SplitCLK_6_339(net1279,net1280_c1,net1281_c1);
SPLITT SplitCLK_6_340(net1268,net1278_c1,net1279_c1);
SPLITT SplitCLK_4_341(net1275,net1276_c1,net1277_c1);
SPLITT SplitCLK_0_342(net1270,net1275_c1,net1274_c1);
SPLITT SplitCLK_6_343(net1271,net1272_c1,net1273_c1);
SPLITT SplitCLK_4_344(net1269,net1271_c1,net1270_c1);
SPLITT SplitCLK_6_345(net1250,net1268_c1,net1269_c1);
SPLITT SplitCLK_0_346(net1265,net1266_c1,net1267_c1);
SPLITT SplitCLK_0_347(net1260,net1265_c1,net1264_c1);
SPLITT SplitCLK_2_348(net1261,net1263_c1,net1262_c1);
SPLITT SplitCLK_6_349(net1252,net1260_c1,net1261_c1);
SPLITT SplitCLK_0_350(net1254,net1259_c1,net1258_c1);
SPLITT SplitCLK_2_351(net1255,net1256_c1,net1257_c1);
SPLITT SplitCLK_4_352(net1253,net1255_c1,net1254_c1);
SPLITT SplitCLK_6_353(net1251,net1253_c1,net1252_c1);
SPLITT SplitCLK_6_354(net1214,net1250_c1,net1251_c1);
SPLITT SplitCLK_4_355(net1247,net1248_c1,net1249_c1);
SPLITT SplitCLK_0_356(net1242,net1247_c1,net1246_c1);
SPLITT SplitCLK_2_357(net1243,net1245_c1,net1244_c1);
SPLITT SplitCLK_4_358(net1234,net1243_c1,net1242_c1);
SPLITT SplitCLK_0_359(net1236,net1241_c1,net1240_c1);
SPLITT SplitCLK_4_360(net1237,net1239_c1,net1238_c1);
SPLITT SplitCLK_4_361(net1235,net1237_c1,net1236_c1);
SPLITT SplitCLK_0_362(net1216,net1234_c1,net1235_c1);
SPLITT SplitCLK_4_363(net1231,net1233_c1,net1232_c1);
SPLITT SplitCLK_4_364(net1226,net1231_c1,net1230_c1);
SPLITT SplitCLK_2_365(net1227,net1228_c1,net1229_c1);
SPLITT SplitCLK_6_366(net1218,net1226_c1,net1227_c1);
SPLITT SplitCLK_4_367(net1220,net1224_c1,net1225_c1);
SPLITT SplitCLK_2_368(net1221,net1222_c1,net1223_c1);
SPLITT SplitCLK_4_369(net1219,net1221_c1,net1220_c1);
SPLITT SplitCLK_4_370(net1217,net1218_c1,net1219_c1);
SPLITT SplitCLK_4_371(net1215,net1217_c1,net1216_c1);
SPLITT SplitCLK_6_372(net1213,net1214_c1,net1215_c1);
SPLITT SplitCLK_6_373(net1062,net1212_c1,net1213_c1);
SPLITT SplitCLK_4_374(net1209,net1210_c1,net1211_c1);
SPLITT SplitCLK_4_375(net1204,net1209_c1,net1208_c1);
SPLITT SplitCLK_6_376(net1205,net1207_c1,net1206_c1);
SPLITT SplitCLK_6_377(net1194,net1204_c1,net1205_c1);
SPLITT SplitCLK_4_378(net1201,net1202_c1,net1203_c1);
SPLITT SplitCLK_0_379(net1196,net1201_c1,net1200_c1);
SPLITT SplitCLK_2_380(net1197,net1199_c1,net1198_c1);
SPLITT SplitCLK_6_381(net1195,net1196_c1,net1197_c1);
SPLITT SplitCLK_4_382(net1176,net1195_c1,net1194_c1);
SPLITT SplitCLK_4_383(net1191,net1192_c1,net1193_c1);
SPLITT SplitCLK_2_384(net1186,net1190_c1,net1191_c1);
SPLITT SplitCLK_6_385(net1187,net1188_c1,net1189_c1);
SPLITT SplitCLK_6_386(net1178,net1186_c1,net1187_c1);
SPLITT SplitCLK_0_387(net1180,net1184_c1,net1185_c1);
SPLITT SplitCLK_4_388(net1181,net1182_c1,net1183_c1);
SPLITT SplitCLK_4_389(net1179,net1181_c1,net1180_c1);
SPLITT SplitCLK_2_390(net1177,net1179_c1,net1178_c1);
SPLITT SplitCLK_6_391(net1138,net1176_c1,net1177_c1);
SPLITT SplitCLK_0_392(net1173,net1174_c1,net1175_c1);
SPLITT SplitCLK_0_393(net1168,net1173_c1,net1172_c1);
SPLITT SplitCLK_6_394(net1169,net1171_c1,net1170_c1);
SPLITT SplitCLK_0_395(net1158,net1169_c1,net1168_c1);
SPLITT SplitCLK_4_396(net1165,net1166_c1,net1167_c1);
SPLITT SplitCLK_4_397(net1160,net1164_c1,net1165_c1);
SPLITT SplitCLK_4_398(net1161,net1163_c1,net1162_c1);
SPLITT SplitCLK_4_399(net1159,net1161_c1,net1160_c1);
SPLITT SplitCLK_0_400(net1140,net1158_c1,net1159_c1);
SPLITT SplitCLK_4_401(net1155,net1156_c1,net1157_c1);
SPLITT SplitCLK_4_402(net1150,net1155_c1,net1154_c1);
SPLITT SplitCLK_6_403(net1151,net1152_c1,net1153_c1);
SPLITT SplitCLK_6_404(net1142,net1150_c1,net1151_c1);
SPLITT SplitCLK_4_405(net1144,net1148_c1,net1149_c1);
SPLITT SplitCLK_6_406(net1145,net1146_c1,net1147_c1);
SPLITT SplitCLK_4_407(net1143,net1145_c1,net1144_c1);
SPLITT SplitCLK_2_408(net1141,net1143_c1,net1142_c1);
SPLITT SplitCLK_4_409(net1139,net1141_c1,net1140_c1);
SPLITT SplitCLK_0_410(net1064,net1138_c1,net1139_c1);
SPLITT SplitCLK_4_411(net1135,net1137_c1,net1136_c1);
SPLITT SplitCLK_4_412(net1130,net1134_c1,net1135_c1);
SPLITT SplitCLK_2_413(net1131,net1132_c1,net1133_c1);
SPLITT SplitCLK_4_414(net1120,net1131_c1,net1130_c1);
SPLITT SplitCLK_4_415(net1127,net1129_c1,net1128_c1);
SPLITT SplitCLK_4_416(net1122,net1127_c1,net1126_c1);
SPLITT SplitCLK_2_417(net1123,net1125_c1,net1124_c1);
SPLITT SplitCLK_4_418(net1121,net1123_c1,net1122_c1);
SPLITT SplitCLK_0_419(net1102,net1120_c1,net1121_c1);
SPLITT SplitCLK_4_420(net1117,net1119_c1,net1118_c1);
SPLITT SplitCLK_0_421(net1112,net1117_c1,net1116_c1);
SPLITT SplitCLK_6_422(net1113,net1115_c1,net1114_c1);
SPLITT SplitCLK_6_423(net1104,net1112_c1,net1113_c1);
SPLITT SplitCLK_0_424(net1106,net1111_c1,net1110_c1);
SPLITT SplitCLK_2_425(net1107,net1109_c1,net1108_c1);
SPLITT SplitCLK_0_426(net1105,net1107_c1,net1106_c1);
SPLITT SplitCLK_2_427(net1103,net1105_c1,net1104_c1);
SPLITT SplitCLK_6_428(net1066,net1102_c1,net1103_c1);
SPLITT SplitCLK_4_429(net1099,net1101_c1,net1100_c1);
SPLITT SplitCLK_0_430(net1094,net1099_c1,net1098_c1);
SPLITT SplitCLK_4_431(net1095,net1096_c1,net1097_c1);
SPLITT SplitCLK_6_432(net1086,net1094_c1,net1095_c1);
SPLITT SplitCLK_4_433(net1088,net1093_c1,net1092_c1);
SPLITT SplitCLK_6_434(net1089,net1090_c1,net1091_c1);
SPLITT SplitCLK_4_435(net1087,net1089_c1,net1088_c1);
SPLITT SplitCLK_0_436(net1068,net1086_c1,net1087_c1);
SPLITT SplitCLK_4_437(net1083,net1084_c1,net1085_c1);
SPLITT SplitCLK_4_438(net1078,net1082_c1,net1083_c1);
SPLITT SplitCLK_6_439(net1079,net1080_c1,net1081_c1);
SPLITT SplitCLK_0_440(net1070,net1079_c1,net1078_c1);
SPLITT SplitCLK_4_441(net1072,net1077_c1,net1076_c1);
SPLITT SplitCLK_2_442(net1073,net1075_c1,net1074_c1);
SPLITT SplitCLK_2_443(net1071,net1072_c1,net1073_c1);
SPLITT SplitCLK_6_444(net1069,net1070_c1,net1071_c1);
SPLITT SplitCLK_4_445(net1067,net1069_c1,net1068_c1);
SPLITT SplitCLK_2_446(net1065,net1067_c1,net1066_c1);
SPLITT SplitCLK_4_447(net1063,net1065_c1,net1064_c1);
SPLITT SplitCLK_0_448(net551,net1062_c1,net1063_c1);
SPLITT SplitCLK_4_449(net1059,net1060_c1,net1061_c1);
SPLITT SplitCLK_4_450(net1054,net1058_c1,net1059_c1);
SPLITT SplitCLK_6_451(net1055,net1056_c1,net1057_c1);
SPLITT SplitCLK_0_452(net1044,net1055_c1,net1054_c1);
SPLITT SplitCLK_4_453(net1051,net1053_c1,net1052_c1);
SPLITT SplitCLK_0_454(net1046,net1051_c1,net1050_c1);
SPLITT SplitCLK_6_455(net1047,net1049_c1,net1048_c1);
SPLITT SplitCLK_4_456(net1045,net1047_c1,net1046_c1);
SPLITT SplitCLK_4_457(net1026,net1044_c1,net1045_c1);
SPLITT SplitCLK_4_458(net1041,net1042_c1,net1043_c1);
SPLITT SplitCLK_0_459(net1036,net1041_c1,net1040_c1);
SPLITT SplitCLK_2_460(net1037,net1039_c1,net1038_c1);
SPLITT SplitCLK_6_461(net1028,net1036_c1,net1037_c1);
SPLITT SplitCLK_4_462(net1030,net1035_c1,net1034_c1);
SPLITT SplitCLK_2_463(net1031,net1033_c1,net1032_c1);
SPLITT SplitCLK_4_464(net1029,net1031_c1,net1030_c1);
SPLITT SplitCLK_6_465(net1027,net1028_c1,net1029_c1);
SPLITT SplitCLK_6_466(net988,net1026_c1,net1027_c1);
SPLITT SplitCLK_4_467(net1023,net1025_c1,net1024_c1);
SPLITT SplitCLK_0_468(net1018,net1023_c1,net1022_c1);
SPLITT SplitCLK_6_469(net1019,net1020_c1,net1021_c1);
SPLITT SplitCLK_6_470(net1008,net1018_c1,net1019_c1);
SPLITT SplitCLK_4_471(net1015,net1017_c1,net1016_c1);
SPLITT SplitCLK_4_472(net1010,net1015_c1,net1014_c1);
SPLITT SplitCLK_2_473(net1011,net1012_c1,net1013_c1);
SPLITT SplitCLK_4_474(net1009,net1011_c1,net1010_c1);
SPLITT SplitCLK_0_475(net990,net1008_c1,net1009_c1);
SPLITT SplitCLK_4_476(net1005,net1006_c1,net1007_c1);
SPLITT SplitCLK_4_477(net1000,net1005_c1,net1004_c1);
SPLITT SplitCLK_6_478(net1001,net1003_c1,net1002_c1);
SPLITT SplitCLK_6_479(net992,net1000_c1,net1001_c1);
SPLITT SplitCLK_0_480(net994,net999_c1,net998_c1);
SPLITT SplitCLK_6_481(net995,net996_c1,net997_c1);
SPLITT SplitCLK_2_482(net993,net994_c1,net995_c1);
SPLITT SplitCLK_2_483(net991,net993_c1,net992_c1);
SPLITT SplitCLK_4_484(net989,net991_c1,net990_c1);
SPLITT SplitCLK_0_485(net914,net988_c1,net989_c1);
SPLITT SplitCLK_4_486(net985,net986_c1,net987_c1);
SPLITT SplitCLK_0_487(net980,net985_c1,net984_c1);
SPLITT SplitCLK_6_488(net981,net982_c1,net983_c1);
SPLITT SplitCLK_6_489(net970,net980_c1,net981_c1);
SPLITT SplitCLK_4_490(net977,net979_c1,net978_c1);
SPLITT SplitCLK_2_491(net972,net976_c1,net977_c1);
SPLITT SplitCLK_6_492(net973,net974_c1,net975_c1);
SPLITT SplitCLK_4_493(net971,net973_c1,net972_c1);
SPLITT SplitCLK_0_494(net952,net970_c1,net971_c1);
SPLITT SplitCLK_0_495(net967,net968_c1,net969_c1);
SPLITT SplitCLK_0_496(net962,net967_c1,net966_c1);
SPLITT SplitCLK_2_497(net963,net964_c1,net965_c1);
SPLITT SplitCLK_0_498(net954,net963_c1,net962_c1);
SPLITT SplitCLK_4_499(net956,net960_c1,net961_c1);
SPLITT SplitCLK_6_500(net957,net958_c1,net959_c1);
SPLITT SplitCLK_4_501(net955,net957_c1,net956_c1);
SPLITT SplitCLK_2_502(net953,net955_c1,net954_c1);
SPLITT SplitCLK_6_503(net916,net952_c1,net953_c1);
SPLITT SplitCLK_4_504(net949,net951_c1,net950_c1);
SPLITT SplitCLK_4_505(net944,net948_c1,net949_c1);
SPLITT SplitCLK_4_506(net945,net946_c1,net947_c1);
SPLITT SplitCLK_6_507(net936,net944_c1,net945_c1);
SPLITT SplitCLK_0_508(net938,net943_c1,net942_c1);
SPLITT SplitCLK_6_509(net939,net941_c1,net940_c1);
SPLITT SplitCLK_4_510(net937,net939_c1,net938_c1);
SPLITT SplitCLK_0_511(net918,net936_c1,net937_c1);
SPLITT SplitCLK_4_512(net933,net934_c1,net935_c1);
SPLITT SplitCLK_4_513(net928,net933_c1,net932_c1);
SPLITT SplitCLK_6_514(net929,net930_c1,net931_c1);
SPLITT SplitCLK_6_515(net920,net928_c1,net929_c1);
SPLITT SplitCLK_4_516(net922,net927_c1,net926_c1);
SPLITT SplitCLK_6_517(net923,net924_c1,net925_c1);
SPLITT SplitCLK_4_518(net921,net923_c1,net922_c1);
SPLITT SplitCLK_4_519(net919,net920_c1,net921_c1);
SPLITT SplitCLK_4_520(net917,net919_c1,net918_c1);
SPLITT SplitCLK_2_521(net915,net917_c1,net916_c1);
SPLITT SplitCLK_6_522(net766,net914_c1,net915_c1);
SPLITT SplitCLK_4_523(net911,net913_c1,net912_c1);
SPLITT SplitCLK_0_524(net906,net911_c1,net910_c1);
SPLITT SplitCLK_6_525(net907,net908_c1,net909_c1);
SPLITT SplitCLK_6_526(net896,net906_c1,net907_c1);
SPLITT SplitCLK_4_527(net903,net904_c1,net905_c1);
SPLITT SplitCLK_0_528(net898,net903_c1,net902_c1);
SPLITT SplitCLK_6_529(net899,net900_c1,net901_c1);
SPLITT SplitCLK_4_530(net897,net899_c1,net898_c1);
SPLITT SplitCLK_0_531(net878,net896_c1,net897_c1);
SPLITT SplitCLK_4_532(net893,net895_c1,net894_c1);
SPLITT SplitCLK_4_533(net888,net893_c1,net892_c1);
SPLITT SplitCLK_0_534(net889,net890_c1,net891_c1);
SPLITT SplitCLK_2_535(net880,net889_c1,net888_c1);
SPLITT SplitCLK_4_536(net882,net887_c1,net886_c1);
SPLITT SplitCLK_2_537(net883,net884_c1,net885_c1);
SPLITT SplitCLK_4_538(net881,net883_c1,net882_c1);
SPLITT SplitCLK_2_539(net879,net881_c1,net880_c1);
SPLITT SplitCLK_6_540(net842,net878_c1,net879_c1);
SPLITT SplitCLK_4_541(net875,net877_c1,net876_c1);
SPLITT SplitCLK_4_542(net870,net875_c1,net874_c1);
SPLITT SplitCLK_2_543(net871,net872_c1,net873_c1);
SPLITT SplitCLK_4_544(net862,net871_c1,net870_c1);
SPLITT SplitCLK_0_545(net864,net868_c1,net869_c1);
SPLITT SplitCLK_4_546(net865,net867_c1,net866_c1);
SPLITT SplitCLK_4_547(net863,net865_c1,net864_c1);
SPLITT SplitCLK_0_548(net844,net862_c1,net863_c1);
SPLITT SplitCLK_4_549(net859,net860_c1,net861_c1);
SPLITT SplitCLK_0_550(net854,net859_c1,net858_c1);
SPLITT SplitCLK_2_551(net855,net857_c1,net856_c1);
SPLITT SplitCLK_6_552(net846,net854_c1,net855_c1);
SPLITT SplitCLK_0_553(net848,net852_c1,net853_c1);
SPLITT SplitCLK_6_554(net849,net850_c1,net851_c1);
SPLITT SplitCLK_4_555(net847,net849_c1,net848_c1);
SPLITT SplitCLK_2_556(net845,net847_c1,net846_c1);
SPLITT SplitCLK_4_557(net843,net845_c1,net844_c1);
SPLITT SplitCLK_6_558(net768,net842_c1,net843_c1);
SPLITT SplitCLK_4_559(net839,net841_c1,net840_c1);
SPLITT SplitCLK_0_560(net834,net839_c1,net838_c1);
SPLITT SplitCLK_6_561(net835,net836_c1,net837_c1);
SPLITT SplitCLK_4_562(net824,net835_c1,net834_c1);
SPLITT SplitCLK_4_563(net831,net833_c1,net832_c1);
SPLITT SplitCLK_4_564(net826,net831_c1,net830_c1);
SPLITT SplitCLK_2_565(net827,net828_c1,net829_c1);
SPLITT SplitCLK_4_566(net825,net827_c1,net826_c1);
SPLITT SplitCLK_0_567(net806,net824_c1,net825_c1);
SPLITT SplitCLK_4_568(net821,net823_c1,net822_c1);
SPLITT SplitCLK_4_569(net816,net821_c1,net820_c1);
SPLITT SplitCLK_6_570(net817,net818_c1,net819_c1);
SPLITT SplitCLK_6_571(net808,net816_c1,net817_c1);
SPLITT SplitCLK_0_572(net810,net815_c1,net814_c1);
SPLITT SplitCLK_0_573(net811,net812_c1,net813_c1);
SPLITT SplitCLK_4_574(net809,net810_c1,net811_c1);
SPLITT SplitCLK_2_575(net807,net809_c1,net808_c1);
SPLITT SplitCLK_6_576(net770,net806_c1,net807_c1);
SPLITT SplitCLK_4_577(net803,net805_c1,net804_c1);
SPLITT SplitCLK_4_578(net798,net802_c1,net803_c1);
SPLITT SplitCLK_6_579(net799,net800_c1,net801_c1);
SPLITT SplitCLK_6_580(net790,net798_c1,net799_c1);
SPLITT SplitCLK_0_581(net792,net796_c1,net797_c1);
SPLITT SplitCLK_2_582(net793,net794_c1,net795_c1);
SPLITT SplitCLK_4_583(net791,net793_c1,net792_c1);
SPLITT SplitCLK_0_584(net772,net790_c1,net791_c1);
SPLITT SplitCLK_4_585(net787,net788_c1,net789_c1);
SPLITT SplitCLK_4_586(net782,net787_c1,net786_c1);
SPLITT SplitCLK_6_587(net783,net784_c1,net785_c1);
SPLITT SplitCLK_6_588(net774,net782_c1,net783_c1);
SPLITT SplitCLK_4_589(net776,net781_c1,net780_c1);
SPLITT SplitCLK_6_590(net777,net778_c1,net779_c1);
SPLITT SplitCLK_4_591(net775,net777_c1,net776_c1);
SPLITT SplitCLK_2_592(net773,net775_c1,net774_c1);
SPLITT SplitCLK_4_593(net771,net773_c1,net772_c1);
SPLITT SplitCLK_2_594(net769,net771_c1,net770_c1);
SPLITT SplitCLK_4_595(net767,net769_c1,net768_c1);
SPLITT SplitCLK_2_596(net552,net767_c1,net766_c1);
wire dummy0;
SPLITT SplitCLK_4_597(net1040,net765_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_4_598(net964,net764_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_599(net796,net763_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_600(net1262,net762_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_601(net1038,net761_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_4_602(net1056,net760_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_2_603(net1182,net759_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_4_604(net1230,net758_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_4_605(net874,net757_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_4_606(net1110,net756_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_2_607(net1132,net755_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_2_608(net1134,net754_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_4_609(net1152,net753_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_2_610(net1188,net752_c1,dummy13);
wire dummy14;
SPLITT SplitCLK_2_611(net1170,net751_c1,dummy14);
wire dummy15;
SPLITT SplitCLK_4_612(net1208,net750_c1,dummy15);
wire dummy16;
SPLITT SplitCLK_4_613(net1332,net749_c1,dummy16);
wire dummy17;
SPLITT SplitCLK_4_614(net1200,net748_c1,dummy17);
wire dummy18;
SPLITT SplitCLK_4_615(net1126,net747_c1,dummy18);
wire dummy19;
SPLITT SplitCLK_4_616(net948,net746_c1,dummy19);
wire dummy20;
SPLITT SplitCLK_4_617(net838,net745_c1,dummy20);
wire dummy21;
SPLITT SplitCLK_2_618(net1153,net744_c1,dummy21);
wire dummy22;
SPLITT SplitCLK_2_619(net1294,net743_c1,dummy22);
wire dummy23;
SPLITT SplitCLK_2_620(net1222,net742_c1,dummy23);
wire dummy24;
SPLITT SplitCLK_2_621(net1224,net741_c1,dummy24);
wire dummy25;
SPLITT SplitCLK_4_622(net1240,net740_c1,dummy25);
wire dummy26;
SPLITT SplitCLK_2_623(net1238,net739_c1,dummy26);
wire dummy27;
SPLITT SplitCLK_2_624(net1296,net738_c1,dummy27);
wire dummy28;
SPLITT SplitCLK_2_625(net974,net737_c1,dummy28);
wire dummy29;
SPLITT SplitCLK_4_626(net1263,net736_c1,dummy29);
wire dummy30;
SPLITT SplitCLK_2_627(net1048,net735_c1,dummy30);
wire dummy31;
SPLITT SplitCLK_2_628(net1300,net734_c1,dummy31);
wire dummy32;
SPLITT SplitCLK_4_629(net1256,net733_c1,dummy32);
wire dummy33;
SPLITT SplitCLK_2_630(net872,net732_c1,dummy33);
wire dummy34;
SPLITT SplitCLK_4_631(net1330,net731_c1,dummy34);
wire dummy35;
SPLITT SplitCLK_4_632(net828,net730_c1,dummy35);
wire dummy36;
SPLITT SplitCLK_4_633(net1111,net729_c1,dummy36);
wire dummy37;
SPLITT SplitCLK_2_634(net1020,net728_c1,dummy37);
wire dummy38;
SPLITT SplitCLK_2_635(net996,net727_c1,dummy38);
wire dummy39;
SPLITT SplitCLK_2_636(net866,net726_c1,dummy39);
wire dummy40;
SPLITT SplitCLK_2_637(net873,net725_c1,dummy40);
wire dummy41;
SPLITT SplitCLK_2_638(net1244,net724_c1,dummy41);
wire dummy42;
SPLITT SplitCLK_4_639(net830,net723_c1,dummy42);
wire dummy43;
SPLITT SplitCLK_2_640(net890,net722_c1,dummy43);
wire dummy44;
SPLITT SplitCLK_4_641(net858,net721_c1,dummy44);
wire dummy45;
SPLITT SplitCLK_2_642(net997,net720_c1,dummy45);
wire dummy46;
SPLITT SplitCLK_4_643(net850,net719_c1,dummy46);
wire dummy47;
SPLITT SplitCLK_2_644(net1114,net718_c1,dummy47);
wire dummy48;
SPLITT SplitCLK_2_645(net778,net717_c1,dummy48);
wire dummy49;
SPLITT SplitCLK_2_646(net1012,net716_c1,dummy49);
wire dummy50;
SPLITT SplitCLK_4_647(net1080,net715_c1,dummy50);
wire dummy51;
SPLITT SplitCLK_2_648(net1223,net714_c1,dummy51);
wire dummy52;
SPLITT SplitCLK_2_649(net1074,net713_c1,dummy52);
wire dummy53;
SPLITT SplitCLK_4_650(net910,net712_c1,dummy53);
wire dummy54;
SPLITT SplitCLK_2_651(net900,net711_c1,dummy54);
wire dummy55;
SPLITT SplitCLK_4_652(net1116,net710_c1,dummy55);
wire dummy56;
SPLITT SplitCLK_4_653(net902,net709_c1,dummy56);
wire dummy57;
SPLITT SplitCLK_4_654(net908,net708_c1,dummy57);
wire dummy58;
SPLITT SplitCLK_2_655(net800,net707_c1,dummy58);
wire dummy59;
SPLITT SplitCLK_4_656(net1098,net706_c1,dummy59);
wire dummy60;
SPLITT SplitCLK_2_657(net856,net705_c1,dummy60);
wire dummy61;
SPLITT SplitCLK_2_658(net901,net704_c1,dummy61);
wire dummy62;
SPLITT SplitCLK_2_659(net836,net703_c1,dummy62);
wire dummy63;
SPLITT SplitCLK_2_660(net1108,net702_c1,dummy63);
wire dummy64;
SPLITT SplitCLK_4_661(net797,net701_c1,dummy64);
wire dummy65;
SPLITT SplitCLK_2_662(net802,net700_c1,dummy65);
wire dummy66;
SPLITT SplitCLK_2_663(net1096,net699_c1,dummy66);
wire dummy67;
SPLITT SplitCLK_2_664(net801,net698_c1,dummy67);
wire dummy68;
SPLITT SplitCLK_2_665(net965,net697_c1,dummy68);
wire dummy69;
SPLITT SplitCLK_4_666(net1050,net696_c1,dummy69);
wire dummy70;
SPLITT SplitCLK_2_667(net946,net695_c1,dummy70);
wire dummy71;
SPLITT SplitCLK_4_668(net942,net694_c1,dummy71);
wire dummy72;
SPLITT SplitCLK_4_669(net1246,net693_c1,dummy72);
wire dummy73;
SPLITT SplitCLK_2_670(net909,net692_c1,dummy73);
wire dummy74;
SPLITT SplitCLK_2_671(net1124,net691_c1,dummy74);
wire dummy75;
SPLITT SplitCLK_4_672(net1258,net690_c1,dummy75);
wire dummy76;
SPLITT SplitCLK_4_673(net1014,net689_c1,dummy76);
wire dummy77;
SPLITT SplitCLK_4_674(net998,net688_c1,dummy77);
wire dummy78;
SPLITT SplitCLK_4_675(net1109,net687_c1,dummy78);
wire dummy79;
SPLITT SplitCLK_4_676(net1115,net686_c1,dummy79);
wire dummy80;
SPLITT SplitCLK_2_677(net1198,net685_c1,dummy80);
wire dummy81;
SPLITT SplitCLK_2_678(net1190,net684_c1,dummy81);
wire dummy82;
SPLITT SplitCLK_4_679(net1310,net683_c1,dummy82);
wire dummy83;
SPLITT SplitCLK_2_680(net1206,net682_c1,dummy83);
wire dummy84;
SPLITT SplitCLK_2_681(net1133,net681_c1,dummy84);
wire dummy85;
SPLITT SplitCLK_4_682(net1320,net680_c1,dummy85);
wire dummy86;
SPLITT SplitCLK_2_683(net1189,net679_c1,dummy86);
wire dummy87;
SPLITT SplitCLK_4_684(net1207,net678_c1,dummy87);
wire dummy88;
SPLITT SplitCLK_2_685(net1311,net677_c1,dummy88);
wire dummy89;
SPLITT SplitCLK_2_686(net1057,net676_c1,dummy89);
wire dummy90;
SPLITT SplitCLK_2_687(net930,net675_c1,dummy90);
wire dummy91;
SPLITT SplitCLK_2_688(net940,net674_c1,dummy91);
wire dummy92;
SPLITT SplitCLK_2_689(net812,net673_c1,dummy92);
wire dummy93;
SPLITT SplitCLK_4_690(net886,net672_c1,dummy93);
wire dummy94;
SPLITT SplitCLK_4_691(net1125,net671_c1,dummy94);
wire dummy95;
SPLITT SplitCLK_4_692(net884,net670_c1,dummy95);
wire dummy96;
SPLITT SplitCLK_2_693(net1239,net669_c1,dummy96);
wire dummy97;
SPLITT SplitCLK_2_694(net887,net668_c1,dummy97);
wire dummy98;
SPLITT SplitCLK_2_695(net1228,net667_c1,dummy98);
wire dummy99;
SPLITT SplitCLK_4_696(net868,net666_c1,dummy99);
wire dummy100;
SPLITT SplitCLK_2_697(net1082,net665_c1,dummy100);
wire dummy101;
SPLITT SplitCLK_4_698(net966,net664_c1,dummy101);
wire dummy102;
SPLITT SplitCLK_4_699(net1146,net663_c1,dummy102);
wire dummy103;
SPLITT SplitCLK_2_700(net867,net662_c1,dummy103);
wire dummy104;
SPLITT SplitCLK_4_701(net794,net661_c1,dummy104);
wire dummy105;
SPLITT SplitCLK_2_702(net1032,net660_c1,dummy105);
wire dummy106;
SPLITT SplitCLK_2_703(net1147,net659_c1,dummy106);
wire dummy107;
SPLITT SplitCLK_4_704(net852,net658_c1,dummy107);
wire dummy108;
SPLITT SplitCLK_4_705(net786,net657_c1,dummy108);
wire dummy109;
SPLITT SplitCLK_2_706(net795,net656_c1,dummy109);
wire dummy110;
SPLITT SplitCLK_4_707(net780,net655_c1,dummy110);
wire dummy111;
SPLITT SplitCLK_4_708(net1154,net654_c1,dummy111);
wire dummy112;
SPLITT SplitCLK_4_709(net818,net653_c1,dummy112);
wire dummy113;
SPLITT SplitCLK_4_710(net958,net652_c1,dummy113);
wire dummy114;
SPLITT SplitCLK_2_711(net781,net651_c1,dummy114);
wire dummy115;
SPLITT SplitCLK_2_712(net1097,net650_c1,dummy115);
wire dummy116;
SPLITT SplitCLK_4_713(net784,net649_c1,dummy116);
wire dummy117;
SPLITT SplitCLK_4_714(net1354,net648_c1,dummy117);
wire dummy118;
SPLITT SplitCLK_4_715(net814,net647_c1,dummy118);
wire dummy119;
SPLITT SplitCLK_2_716(net924,net646_c1,dummy119);
wire dummy120;
SPLITT SplitCLK_2_717(net1081,net645_c1,dummy120);
wire dummy121;
SPLITT SplitCLK_4_718(net820,net644_c1,dummy121);
wire dummy122;
SPLITT SplitCLK_4_719(net1280,net643_c1,dummy122);
wire dummy123;
SPLITT SplitCLK_2_720(net819,net642_c1,dummy123);
wire dummy124;
SPLITT SplitCLK_2_721(net960,net641_c1,dummy124);
wire dummy125;
SPLITT SplitCLK_4_722(net779,net640_c1,dummy125);
wire dummy126;
SPLITT SplitCLK_4_723(net941,net639_c1,dummy126);
wire dummy127;
SPLITT SplitCLK_4_724(net926,net638_c1,dummy127);
wire dummy128;
SPLITT SplitCLK_4_725(net932,net637_c1,dummy128);
wire dummy129;
SPLITT SplitCLK_2_726(net829,net636_c1,dummy129);
wire dummy130;
SPLITT SplitCLK_2_727(net1281,net635_c1,dummy130);
wire dummy131;
SPLITT SplitCLK_4_728(net925,net634_c1,dummy131);
wire dummy132;
SPLITT SplitCLK_4_729(net961,net633_c1,dummy132);
wire dummy133;
SPLITT SplitCLK_4_730(net1022,net632_c1,dummy133);
wire dummy134;
SPLITT SplitCLK_2_731(net1257,net631_c1,dummy134);
wire dummy135;
SPLITT SplitCLK_4_732(net1295,net630_c1,dummy135);
wire dummy136;
SPLITT SplitCLK_4_733(net1297,net629_c1,dummy136);
wire dummy137;
SPLITT SplitCLK_4_734(net1092,net628_c1,dummy137);
wire dummy138;
SPLITT SplitCLK_2_735(net1331,net627_c1,dummy138);
wire dummy139;
SPLITT SplitCLK_2_736(net927,net626_c1,dummy139);
wire dummy140;
SPLITT SplitCLK_4_737(net975,net625_c1,dummy140);
wire dummy141;
SPLITT SplitCLK_2_738(net1164,net624_c1,dummy141);
wire dummy142;
SPLITT SplitCLK_2_739(net1002,net623_c1,dummy142);
wire dummy143;
SPLITT SplitCLK_4_740(net1336,net622_c1,dummy143);
wire dummy144;
SPLITT SplitCLK_2_741(net976,net621_c1,dummy144);
wire dummy145;
SPLITT SplitCLK_4_742(net1003,net620_c1,dummy145);
wire dummy146;
SPLITT SplitCLK_4_743(net1171,net619_c1,dummy146);
wire dummy147;
SPLITT SplitCLK_4_744(net1199,net618_c1,dummy147);
wire dummy148;
SPLITT SplitCLK_2_745(net1346,net617_c1,dummy148);
wire dummy149;
SPLITT SplitCLK_4_746(net1264,net616_c1,dummy149);
wire dummy150;
SPLITT SplitCLK_4_747(net1049,net615_c1,dummy150);
wire dummy151;
SPLITT SplitCLK_4_748(net1318,net614_c1,dummy151);
wire dummy152;
SPLITT SplitCLK_2_749(net1319,net613_c1,dummy152);
wire dummy153;
SPLITT SplitCLK_4_750(net984,net612_c1,dummy153);
wire dummy154;
SPLITT SplitCLK_4_751(net1034,net611_c1,dummy154);
wire dummy155;
SPLITT SplitCLK_2_752(net815,net610_c1,dummy155);
wire dummy156;
SPLITT SplitCLK_4_753(net1241,net609_c1,dummy156);
wire dummy157;
SPLITT SplitCLK_2_754(net1184,net608_c1,dummy157);
wire dummy158;
SPLITT SplitCLK_4_755(net1162,net607_c1,dummy158);
wire dummy159;
SPLITT SplitCLK_4_756(net891,net606_c1,dummy159);
wire dummy160;
SPLITT SplitCLK_2_757(net1035,net605_c1,dummy160);
wire dummy161;
SPLITT SplitCLK_4_758(net931,net604_c1,dummy161);
wire dummy162;
SPLITT SplitCLK_4_759(net1356,net603_c1,dummy162);
wire dummy163;
SPLITT SplitCLK_2_760(net837,net602_c1,dummy163);
wire dummy164;
SPLITT SplitCLK_2_761(net1093,net601_c1,dummy164);
wire dummy165;
SPLITT SplitCLK_2_762(net1229,net600_c1,dummy165);
wire dummy166;
SPLITT SplitCLK_4_763(net1004,net599_c1,dummy166);
wire dummy167;
SPLITT SplitCLK_2_764(net1301,net598_c1,dummy167);
wire dummy168;
SPLITT SplitCLK_4_765(net1033,net597_c1,dummy168);
wire dummy169;
SPLITT SplitCLK_4_766(net1333,net596_c1,dummy169);
wire dummy170;
SPLITT SplitCLK_2_767(net947,net595_c1,dummy170);
wire dummy171;
SPLITT SplitCLK_4_768(net1347,net594_c1,dummy171);
wire dummy172;
SPLITT SplitCLK_2_769(net1148,net593_c1,dummy172);
wire dummy173;
SPLITT SplitCLK_4_770(net869,net592_c1,dummy173);
wire dummy174;
SPLITT SplitCLK_4_771(net1075,net591_c1,dummy174);
wire dummy175;
SPLITT SplitCLK_4_772(net1348,net590_c1,dummy175);
wire dummy176;
SPLITT SplitCLK_4_773(net892,net589_c1,dummy176);
wire dummy177;
SPLITT SplitCLK_2_774(net1058,net588_c1,dummy177);
wire dummy178;
SPLITT SplitCLK_2_775(net959,net587_c1,dummy178);
wire dummy179;
SPLITT SplitCLK_4_776(net1090,net586_c1,dummy179);
wire dummy180;
SPLITT SplitCLK_2_777(net1013,net585_c1,dummy180);
wire dummy181;
SPLITT SplitCLK_4_778(net1172,net584_c1,dummy181);
wire dummy182;
SPLITT SplitCLK_4_779(net1274,net583_c1,dummy182);
wire dummy183;
SPLITT SplitCLK_4_780(net1338,net582_c1,dummy183);
wire dummy184;
SPLITT SplitCLK_4_781(net982,net581_c1,dummy184);
wire dummy185;
SPLITT SplitCLK_2_782(net1091,net580_c1,dummy185);
wire dummy186;
SPLITT SplitCLK_4_783(net1245,net579_c1,dummy186);
wire dummy187;
SPLITT SplitCLK_4_784(net1076,net578_c1,dummy187);
wire dummy188;
SPLITT SplitCLK_4_785(net999,net577_c1,dummy188);
wire dummy189;
SPLITT SplitCLK_4_786(net813,net576_c1,dummy189);
wire dummy190;
SPLITT SplitCLK_2_787(net1355,net575_c1,dummy190);
wire dummy191;
SPLITT SplitCLK_2_788(net983,net574_c1,dummy191);
wire dummy192;
SPLITT SplitCLK_2_789(net1077,net573_c1,dummy192);
wire dummy193;
SPLITT SplitCLK_2_790(net1312,net572_c1,dummy193);
wire dummy194;
SPLITT SplitCLK_4_791(net1185,net571_c1,dummy194);
wire dummy195;
SPLITT SplitCLK_4_792(net853,net570_c1,dummy195);
wire dummy196;
SPLITT SplitCLK_2_793(net885,net569_c1,dummy196);
wire dummy197;
SPLITT SplitCLK_2_794(net1272,net568_c1,dummy197);
wire dummy198;
SPLITT SplitCLK_4_795(net943,net567_c1,dummy198);
wire dummy199;
SPLITT SplitCLK_4_796(net1302,net566_c1,dummy199);
wire dummy200;
SPLITT SplitCLK_4_797(net1149,net565_c1,dummy200);
wire dummy201;
SPLITT SplitCLK_2_798(net785,net564_c1,dummy201);
wire dummy202;
SPLITT SplitCLK_4_799(net1183,net563_c1,dummy202);
wire dummy203;
SPLITT SplitCLK_2_800(net1259,net562_c1,dummy203);
wire dummy204;
SPLITT SplitCLK_2_801(net1273,net561_c1,dummy204);
wire dummy205;
SPLITT SplitCLK_4_802(net1225,net560_c1,dummy205);
wire dummy206;
SPLITT SplitCLK_2_803(net1163,net559_c1,dummy206);
wire dummy207;
SPLITT SplitCLK_4_804(net857,net558_c1,dummy207);
wire dummy208;
SPLITT SplitCLK_2_805(net1337,net557_c1,dummy208);
wire dummy209;
SPLITT SplitCLK_4_806(net1282,net556_c1,dummy209);
wire dummy210;
SPLITT SplitCLK_4_807(net1039,net555_c1,dummy210);
wire dummy211;
SPLITT SplitCLK_2_808(net1021,net554_c1,dummy211);
wire dummy212;
SPLITT SplitCLK_2_809(net851,net553_c1,dummy212);
SPLITT SplitCLK_0_810(net1360,net551_c1,net552_c1);
wire dummy213;
SPLITT Split_HOLD_943(net408,dummy213,net1361_c1);
wire dummy214;
SPLITT Split_HOLD_944(net399,dummy214,net1362_c1);
wire dummy215;
SPLITT Split_HOLD_945(net506,dummy215,net1363_c1);
INTERCONNECT TMS_Pad_Split_307_n763(TMS_Pad,net0);
INTERCONNECT AND2T_16_n40_Split_317_n773(net1_c1,net1);
INTERCONNECT NOTT_8_n32_Split_311_n767(net2_c1,net2);
INTERCONNECT NOTT_17_n41_AND2T_144_n180(net3_c1,net3);
INTERCONNECT AND2T_9_n33_DFFT_155__PIPL_n209(net4_c1,net4);
INTERCONNECT AND2T_26_n50_Split_328_n784(net5_c1,net5);
INTERCONNECT AND2T_18_n42_Split_318_n774(net6_c1,net6);
INTERCONNECT AND2T_10_n34_DFFT_156__PIPL_n210(net7_c1,net7);
INTERCONNECT AND2T_27_n51_Split_329_n785(net8_c1,net8);
INTERCONNECT NOTT_19_n43_OR2T_100_n124(net9_c1,net9);
INTERCONNECT AND2T_11_n35_DFFT_157__PIPL_n211(net10_c1,net10);
INTERCONNECT XOR2T_36_n60_DFFT_188__FPB_n644(net11_c1,net11);
INTERCONNECT AND2T_28_n52_Split_331_n787(net12_c1,net12);
INTERCONNECT NOTT_20_n44_AND2T_143_n179(net13_c1,net13);
INTERCONNECT AND2T_12_n36_DFFT_158__PIPL_n212(net14_c1,net14);
INTERCONNECT OR2T_37_n61_OR2T_38_n62(net15_c1,net15);
INTERCONNECT AND2T_29_n53_Split_332_n788(net16_c1,net16);
INTERCONNECT AND2T_21_n45_AND2T_114_n138(net17_c1,net17);
INTERCONNECT AND2T_13_n37_DFFT_263__FPB_n719(net18_c1,net18);
INTERCONNECT AND2T_46_n70_DFFT_194__FPB_n650(net19_c1,net19);
INTERCONNECT OR2T_38_n62_NOTT_49_n73(net20_c1,net20);
INTERCONNECT OR2T_30_n54_OR2T_31_n55(net21_c1,net21);
INTERCONNECT AND2T_22_n46_Split_321_n777(net22_c1,net22);
INTERCONNECT NOTT_14_n38_Split_314_n770(net23_c1,net23);
INTERCONNECT NOTT_47_n71_AND2T_46_n70(net24_c1,net24);
INTERCONNECT AND2T_39_n63_Split_336_n792(net25_c1,net25);
INTERCONNECT OR2T_31_n55_OR2T_38_n62(net26_c1,net26);
INTERCONNECT OR2T_23_n47_OR2T_31_n55(net27_c1,net27);
INTERCONNECT AND2T_15_n39_AND2T_114_n138(net28_c1,net28);
INTERCONNECT AND2T_56_n80_OR2T_59_n83(net29_c1,net29);
INTERCONNECT AND2T_48_n72_Split_339_n795(net30_c1,net30);
INTERCONNECT NOTT_40_n64_AND2T_43_n67(net31_c1,net31);
INTERCONNECT AND2T_32_n56_Split_333_n789(net32_c1,net32);
INTERCONNECT AND2T_24_n48_Split_323_n779(net33_c1,net33);
INTERCONNECT AND2T_57_n81_OR2T_59_n83(net34_c1,net34);
INTERCONNECT NOTT_49_n73_AND2T_48_n72(net35_c1,net35);
INTERCONNECT NOTT_41_n65_Split_337_n793(net36_c1,net36);
INTERCONNECT AND2T_33_n57_Split_334_n790(net37_c1,net37);
INTERCONNECT AND2T_25_n49_Split_325_n781(net38_c1,net38);
INTERCONNECT AND2T_66_n90_Split_347_n803(net39_c1,net39);
INTERCONNECT OR2T_58_n82_DFFT_202__FPB_n658(net40_c1,net40);
INTERCONNECT NOTT_50_n74_Split_342_n798(net41_c1,net41);
INTERCONNECT OR2T_42_n66_DFFT_190__FPB_n646(net42_c1,net42);
INTERCONNECT OR2T_34_n58_OR2T_37_n61(net43_c1,net43);
INTERCONNECT AND2T_67_n91_AND2T_68_n92(net44_c1,net44);
INTERCONNECT OR2T_59_n83_OR2T_60_n84(net45_c1,net45);
INTERCONNECT AND2T_51_n75_Split_343_n799(net46_c1,net46);
INTERCONNECT AND2T_43_n67_Split_338_n794(net47_c1,net47);
INTERCONNECT AND2T_35_n59_DFFT_189__FPB_n645(net48_c1,net48);
INTERCONNECT AND2T_68_n92_OR2T_69_n93(net49_c1,net49);
INTERCONNECT OR2T_60_n84_DFFT_214__FPB_n670(net50_c1,net50);
INTERCONNECT AND2T_52_n76_AND2T_53_n77(net51_c1,net51);
INTERCONNECT AND2T_44_n68_NOTT_47_n71(net52_c1,net52);
INTERCONNECT OR2T_69_n93_OR2T_70_n94(net53_c1,net53);
INTERCONNECT AND2T_61_n85_DFFT_205__FPB_n661(net54_c1,net54);
INTERCONNECT AND2T_53_n77_DFFT_204__FPB_n660(net55_c1,net55);
INTERCONNECT XOR2T_45_n69_AND2T_44_n68(net56_c1,net56);
INTERCONNECT OR2T_70_n94_OR2T_75_n99(net57_c1,net57);
INTERCONNECT OR2T_62_n86_AND2T_63_n87(net58_c1,net58);
INTERCONNECT AND2T_54_n78_Split_345_n801(net59_c1,net59);
INTERCONNECT AND2T_71_n95_Split_348_n804(net60_c1,net60);
INTERCONNECT AND2T_63_n87_DFFT_213__FPB_n669(net61_c1,net61);
INTERCONNECT XOR2T_55_n79_DFFT_201__FPB_n657(net62_c1,net62);
INTERCONNECT AND2T_72_n96_OR2T_74_n98(net63_c1,net63);
INTERCONNECT AND2T_64_n88_Split_346_n802(net64_c1,net64);
INTERCONNECT AND2T_73_n97_OR2T_74_n98(net65_c1,net65);
INTERCONNECT OR2T_65_n89_OR2T_70_n94(net66_c1,net66);
INTERCONNECT OR2T_74_n98_OR2T_75_n99(net67_c1,net67);
INTERCONNECT OR2T_75_n99_OR2T_76_n100(net68_c1,net68);
INTERCONNECT OR2T_76_n100_OR2T_77_n101(net69_c1,net69);
INTERCONNECT OR2T_77_n101_OR2T_78_n102(net70_c1,net70);
INTERCONNECT AND2T_86_n110_OR2T_88_n112(net71_c1,net71);
INTERCONNECT OR2T_78_n102_AND2T_80_n104(net72_c1,net72);
INTERCONNECT AND2T_87_n111_OR2T_88_n112(net73_c1,net73);
INTERCONNECT NOTT_79_n103_DFFT_215__FPB_n671(net74_c1,net74);
INTERCONNECT OR2T_96_n120_AND2T_98_n122(net75_c1,net75);
INTERCONNECT OR2T_88_n112_OR2T_89_n113(net76_c1,net76);
INTERCONNECT AND2T_80_n104_Split_349_n805(net77_c1,net77);
INTERCONNECT NOTT_97_n121_DFFT_233__FPB_n689(net78_c1,net78);
INTERCONNECT OR2T_89_n113_OR2T_94_n118(net79_c1,net79);
INTERCONNECT AND2T_81_n105_OR2T_95_n119(net80_c1,net80);
INTERCONNECT AND2T_106_n130_OR2T_107_n131(net81_c1,net81);
INTERCONNECT AND2T_98_n122_Split_352_n808(net82_c1,net82);
INTERCONNECT AND2T_90_n114_DFFT_229__FPB_n685(net83_c1,net83);
INTERCONNECT NOTT_82_n106_AND2T_81_n105(net84_c1,net84);
INTERCONNECT OR2T_107_n131_OR2T_108_n132(net85_c1,net85);
INTERCONNECT AND2T_99_n123_Split_355_n811(net86_c1,net86);
INTERCONNECT AND2T_91_n115_OR2T_93_n117(net87_c1,net87);
INTERCONNECT AND2T_83_n107_DFFT_227__FPB_n683(net88_c1,net88);
INTERCONNECT OR2T_116_n140_OR2T_117_n141(net89_c1,net89);
INTERCONNECT OR2T_108_n132_OR2T_118_n142(net90_c1,net90);
INTERCONNECT OR2T_100_n124_AND2T_99_n123(net91_c1,net91);
INTERCONNECT AND2T_92_n116_Split_351_n807(net92_c1,net92);
INTERCONNECT AND2T_84_n108_AND2T_83_n107(net93_c1,net93);
INTERCONNECT OR2T_117_n141_OR2T_118_n142(net94_c1,net94);
INTERCONNECT AND2T_109_n133_DFFT_248__FPB_n704(net95_c1,net95);
INTERCONNECT AND2T_101_n125_Split_356_n812(net96_c1,net96);
INTERCONNECT OR2T_93_n117_OR2T_94_n118(net97_c1,net97);
INTERCONNECT AND2T_85_n109_AND2T_86_n110(net98_c1,net98);
INTERCONNECT OR2T_126_n150_OR2T_136_n160(net99_c1,net99);
INTERCONNECT OR2T_118_n142_DFFT_249__FPB_n705(net100_c1,net100);
INTERCONNECT AND2T_110_n134_OR2T_111_n135(net101_c1,net101);
INTERCONNECT OR2T_102_n126_AND2T_103_n127(net102_c1,net102);
INTERCONNECT OR2T_94_n118_DFFT_232__FPB_n688(net103_c1,net103);
INTERCONNECT OR2T_127_n151_AND2T_129_n153(net104_c1,net104);
INTERCONNECT OR2T_119_n143_AND2T_121_n145(net105_c1,net105);
INTERCONNECT OR2T_111_n135_OR2T_112_n136(net106_c1,net106);
INTERCONNECT AND2T_103_n127_DFFT_246__FPB_n702(net107_c1,net107);
INTERCONNECT OR2T_95_n119_OR2T_96_n120(net108_c1,net108);
INTERCONNECT OR2T_136_n160_DFFT_267__FPB_n723(net109_c1,net109);
INTERCONNECT AND2T_128_n152_AND2T_129_n153(net110_c1,net110);
INTERCONNECT NOTT_120_n144_DFFT_250__FPB_n706(net111_c1,net111);
INTERCONNECT OR2T_112_n136_OR2T_117_n141(net112_c1,net112);
INTERCONNECT AND2T_104_n128_OR2T_107_n131(net113_c1,net113);
INTERCONNECT OR2T_137_n161_AND2T_139_n163(net114_c1,net114);
INTERCONNECT AND2T_129_n153_OR2T_131_n155(net115_c1,net115);
INTERCONNECT AND2T_121_n145_Split_360_n816(net116_c1,net116);
INTERCONNECT AND2T_113_n137_Split_358_n814(net117_c1,net117);
INTERCONNECT AND2T_105_n129_Split_357_n813(net118_c1,net118);
INTERCONNECT NOTT_138_n162_DFFT_268__FPB_n724(net119_c1,net119);
INTERCONNECT OR2T_130_n154_OR2T_131_n155(net120_c1,net120);
INTERCONNECT AND2T_122_n146_DFFT_262__FPB_n718(net121_c1,net121);
INTERCONNECT AND2T_114_n138_Split_359_n815(net122_c1,net122);
INTERCONNECT AND2T_139_n163_Split_363_n819(net123_c1,net123);
INTERCONNECT OR2T_131_n155_OR2T_135_n159(net124_c1,net124);
INTERCONNECT AND2T_123_n147_DFFT_261__FPB_n717(net125_c1,net125);
INTERCONNECT OR2T_115_n139_OR2T_116_n140(net126_c1,net126);
INTERCONNECT AND2T_144_n180_Split_375_n831(net127_c1,net127);
INTERCONNECT AND2T_132_n156_OR2T_134_n158(net128_c1,net128);
INTERCONNECT AND2T_124_n148_OR2T_126_n150(net129_c1,net129);
INTERCONNECT AND2T_145_n181_Split_378_n834(net130_c1,net130);
INTERCONNECT AND2T_133_n157_OR2T_134_n158(net131_c1,net131);
INTERCONNECT OR2T_125_n149_AND2T_124_n148(net132_c1,net132);
INTERCONNECT AND2T_146_n182_Split_381_n837(net133_c1,net133);
INTERCONNECT OR2T_134_n158_OR2T_135_n159(net134_c1,net134);
INTERCONNECT NOTT_147_n183_Split_384_n840(net135_c1,net135);
INTERCONNECT OR2T_135_n159_OR2T_136_n160(net136_c1,net136);
INTERCONNECT NOTT_148_n184_Split_387_n843(net137_c1,net137);
INTERCONNECT AND2T_140_n176_Split_365_n821(net138_c1,net138);
INTERCONNECT AND2T_141_n177_Split_368_n824(net139_c1,net139);
INTERCONNECT NOTT_142_n178_Split_371_n827(net140_c1,net140);
INTERCONNECT AND2T_143_n179_Split_372_n828(net141_c1,net141);
INTERCONNECT NOTT_149_n197_Split_390_n846(net142_c1,net142);
INTERCONNECT NOTT_150_n198_Split_393_n849(net143_c1,net143);
INTERCONNECT NOTT_151_n199_Split_396_n852(net144_c1,net144);
INTERCONNECT Split_344_n800_DFFT_197__FPB_n653(net145_c1,net145);
INTERCONNECT Split_345_n801_AND2T_91_n115(net146_c1,net146);
INTERCONNECT Split_354_n810_DFFT_171__FBL_n627(net147_c1,net147);
INTERCONNECT Split_346_n802_OR2T_111_n135(net148_c1,net148);
INTERCONNECT TRST_Pad_Split_310_n766(TRST_Pad,net149);
INTERCONNECT Split_355_n811_OR2T_130_n154(net150_c1,net150);
INTERCONNECT Split_347_n803_AND2T_122_n146(net151_c1,net151);
INTERCONNECT Split_364_n820_DFFT_166__FBL_n622(net152_c1,net152);
INTERCONNECT Split_356_n812_AND2T_110_n134(net153_c1,net153);
INTERCONNECT Split_348_n804_OR2T_130_n154(net154_c1,net154);
INTERCONNECT Split_365_n821_Split_367_n823(net155_c1,net155);
INTERCONNECT Split_349_n805_Split_350_n806(net156_c1,net156);
INTERCONNECT Split_357_n813_DFFT_245__FPB_n701(net157_c1,net157);
INTERCONNECT Split_350_n806_DFFT_163__FBL_n619(net158_c1,net158);
INTERCONNECT Split_358_n814_OR2T_125_n149(net159_c1,net159);
INTERCONNECT Split_366_n822_DFFT_182__FPB_n638(net160_c1,net160);
INTERCONNECT Split_374_n830_AND2T_64_n88(net161_c1,net161);
INTERCONNECT Split_375_n831_Split_377_n833(net162_c1,net162);
INTERCONNECT Split_367_n823_DFFT_247__FPB_n703(net163_c1,net163);
INTERCONNECT Split_359_n815_OR2T_125_n149(net164_c1,net164);
INTERCONNECT Split_351_n807_OR2T_116_n140(net165_c1,net165);
INTERCONNECT Split_384_n840_Split_386_n842(net166_c1,net166);
INTERCONNECT Split_368_n824_Split_370_n826(net167_c1,net167);
INTERCONNECT Split_360_n816_Split_362_n818(net168_c1,net168);
INTERCONNECT Split_352_n808_Split_354_n810(net169_c1,net169);
INTERCONNECT Split_376_n832_AND2T_32_n56(net170_c1,net170);
INTERCONNECT Split_361_n817_DFFT_165__FBL_n621(net171_c1,net171);
INTERCONNECT Split_353_n809_DFFT_164__FBL_n620(net172_c1,net172);
INTERCONNECT Split_385_n841_XOR2T_55_n79(net173_c1,net173);
INTERCONNECT Split_377_n833_AND2T_71_n95(net174_c1,net174);
INTERCONNECT Split_369_n825_AND2T_33_n57(net175_c1,net175);
INTERCONNECT Split_378_n834_Split_380_n836(net176_c1,net176);
INTERCONNECT Split_314_n770_Split_316_n772(net177_c1,net177);
INTERCONNECT Split_362_n818_DFFT_172__FBL_n628(net178_c1,net178);
INTERCONNECT Split_370_n826_AND2T_113_n137(net179_c1,net179);
INTERCONNECT Split_386_n842_DFFT_206__FPB_n662(net180_c1,net180);
INTERCONNECT Split_394_n850_AND2T_24_n48(net181_c1,net181);
INTERCONNECT Split_387_n843_Split_389_n845(net182_c1,net182);
INTERCONNECT Split_307_n763_Split_309_n765(net183_c1,net183);
INTERCONNECT Split_363_n819_Split_364_n820(net184_c1,net184);
INTERCONNECT Split_371_n827_AND2T_145_n181(net185_c1,net185);
INTERCONNECT Split_395_n851_DFFT_193__FPB_n649(net186_c1,net186);
INTERCONNECT Split_379_n835_AND2T_35_n59(net187_c1,net187);
INTERCONNECT Split_315_n771_AND2T_18_n42(net188_c1,net188);
INTERCONNECT Split_396_n852_Split_398_n854(net189_c1,net189);
INTERCONNECT Split_372_n828_Split_374_n830(net190_c1,net190);
INTERCONNECT Split_404_n860_DFFT_265__FPB_n721(net191_c1,net191);
INTERCONNECT Split_308_n764_NOTT_148_n184(net192_c1,net192);
INTERCONNECT Split_316_n772_DFFT_191__FPB_n647(net193_c1,net193);
INTERCONNECT Split_324_n780_AND2T_110_n134(net194_c1,net194);
INTERCONNECT Split_388_n844_DFFT_210__FPB_n666(net195_c1,net195);
INTERCONNECT Split_380_n836_AND2T_66_n90(net196_c1,net196);
INTERCONNECT Split_405_n861_Split_407_n863(net197_c1,net197);
INTERCONNECT Split_381_n837_Split_383_n839(net198_c1,net198);
INTERCONNECT Split_325_n781_Split_327_n783(net199_c1,net199);
INTERCONNECT Split_389_n845_DFFT_242__FPB_n698(net200_c1,net200);
INTERCONNECT Split_309_n765_DFFT_153__FPB_n207(net201_c1,net201);
INTERCONNECT Split_317_n773_AND2T_104_n128(net202_c1,net202);
INTERCONNECT Split_373_n829_AND2T_39_n63(net203_c1,net203);
INTERCONNECT Split_397_n853_AND2T_25_n49(net204_c1,net204);
INTERCONNECT Split_390_n846_Split_392_n848(net205_c1,net205);
INTERCONNECT Split_318_n774_Split_320_n776(net206_c1,net206);
INTERCONNECT Split_310_n766_DFFT_154__FPB_n208(net207_c1,net207);
INTERCONNECT Split_334_n790_Split_335_n791(net208_c1,net208);
INTERCONNECT Split_398_n854_OR2T_100_n124(net209_c1,net209);
INTERCONNECT Split_382_n838_AND2T_61_n85(net210_c1,net210);
INTERCONNECT Split_414_n870_DFFT_259__FPB_n715(net211_c1,net211);
INTERCONNECT Split_326_n782_AND2T_33_n57(net212_c1,net212);
INTERCONNECT Split_406_n862_NOTT_79_n103(net213_c1,net213);
INTERCONNECT Split_399_n855_Split_401_n857(net214_c1,net214);
INTERCONNECT Split_311_n767_Split_313_n769(net215_c1,net215);
INTERCONNECT Split_383_n839_DFFT_196__FPB_n652(net216_c1,net216);
INTERCONNECT Split_415_n871_Split_416_n872(net217_c1,net217);
INTERCONNECT Split_407_n863_NOTT_120_n144(net218_c1,net218);
INTERCONNECT Split_327_n783_OR2T_102_n126(net219_c1,net219);
INTERCONNECT Split_335_n791_AND2T_92_n116(net220_c1,net220);
INTERCONNECT Split_319_n775_AND2T_54_n78(net221_c1,net221);
INTERCONNECT Split_391_n847_AND2T_27_n51(net222_c1,net222);
INTERCONNECT Split_408_n864_Split_409_n865(net223_c1,net223);
INTERCONNECT Split_416_n872_NOTT_142_n178(net224_c1,net224);
INTERCONNECT Split_392_n848_AND2T_83_n107(net225_c1,net225);
INTERCONNECT Split_320_n776_AND2T_109_n133(net226_c1,net226);
INTERCONNECT Split_400_n856_AND2T_67_n91(net227_c1,net227);
INTERCONNECT Split_336_n792_OR2T_62_n86(net228_c1,net228);
INTERCONNECT Split_328_n784_AND2T_132_n156(net229_c1,net229);
INTERCONNECT Split_424_n880_AND2T_28_n52(net230_c1,net230);
INTERCONNECT Split_312_n768_AND2T_10_n34(net231_c1,net231);
INTERCONNECT Split_393_n849_Split_395_n851(net232_c1,net232);
INTERCONNECT Split_409_n865_DFFT_198__FPB_n654(net233_c1,net233);
INTERCONNECT Split_425_n881_DFFT_183__FPB_n639(net234_c1,net234);
INTERCONNECT Split_417_n873_DFFT_278__FPB_n734(net235_c1,net235);
INTERCONNECT Split_329_n785_Split_330_n786(net236_c1,net236);
INTERCONNECT Split_321_n777_Split_322_n778(net237_c1,net237);
INTERCONNECT Split_401_n857_DFFT_222__FPB_n678(net238_c1,net238);
INTERCONNECT Split_337_n793_AND2T_128_n152(net239_c1,net239);
INTERCONNECT Split_313_n769_AND2T_12_n36(net240_c1,net240);
INTERCONNECT Split_426_n882_Split_428_n884(net241_c1,net241);
INTERCONNECT Split_402_n858_Split_404_n860(net242_c1,net242);
INTERCONNECT Split_410_n866_Split_411_n867(net243_c1,net243);
INTERCONNECT Split_418_n874_DFFT_276__FPB_n732(net244_c1,net244);
INTERCONNECT Split_330_n786_AND2T_86_n110(net245_c1,net245);
INTERCONNECT Split_338_n794_NOTT_82_n106(net246_c1,net246);
INTERCONNECT Split_322_n778_AND2T_57_n81(net247_c1,net247);
INTERCONNECT Split_339_n795_Split_341_n797(net248_c1,net248);
INTERCONNECT Split_331_n787_DFFT_240__FPB_n696(net249_c1,net249);
INTERCONNECT Split_419_n875_DFFT_277__FPB_n733(net250_c1,net250);
INTERCONNECT Split_323_n779_Split_324_n780(net251_c1,net251);
INTERCONNECT Split_403_n859_AND2T_105_n129(net252_c1,net252);
INTERCONNECT Split_411_n867_DFFT_200__FPB_n656(net253_c1,net253);
INTERCONNECT Split_427_n883_NOTT_20_n44(net254_c1,net254);
INTERCONNECT Split_420_n876_Split_422_n878(net255_c1,net255);
INTERCONNECT Split_412_n868_Split_413_n869(net256_c1,net256);
INTERCONNECT Split_428_n884_DFFT_185__FPB_n641(net257_c1,net257);
INTERCONNECT Split_340_n796_OR2T_96_n120(net258_c1,net258);
INTERCONNECT Split_332_n788_OR2T_65_n89(net259_c1,net259);
INTERCONNECT Split_429_n885_Split_431_n887(net260_c1,net260);
INTERCONNECT Split_341_n797_OR2T_137_n161(net261_c1,net261);
INTERCONNECT Split_413_n869_AND2T_84_n108(net262_c1,net262);
INTERCONNECT Split_333_n789_AND2T_73_n97(net263_c1,net263);
INTERCONNECT Split_421_n877_NOTT_19_n43(net264_c1,net264);
INTERCONNECT Split_422_n878_DFFT_184__FPB_n640(net265_c1,net265);
INTERCONNECT Split_342_n798_DFFT_264__FPB_n720(net266_c1,net266);
INTERCONNECT Split_430_n886_AND2T_28_n52(net267_c1,net267);
INTERCONNECT Split_423_n879_Split_425_n881(net268_c1,net268);
INTERCONNECT Split_343_n799_Split_344_n800(net269_c1,net269);
INTERCONNECT Split_431_n887_DFFT_181__FPB_n637(net270_c1,net270);
INTERCONNECT Split_344_n800_AND2T_87_n111(net271_c1,net271);
INTERCONNECT Split_345_n801_AND2T_56_n80(net272_c1,net272);
INTERCONNECT Split_346_n802_OR2T_65_n89(net273_c1,net273);
INTERCONNECT Split_354_n810_DFFT_168__FBL_n624(net274_c1,net274);
INTERCONNECT Split_347_n803_OR2T_69_n93(net275_c1,net275);
INTERCONNECT Split_355_n811_AND2T_103_n127(net276_c1,net276);
INTERCONNECT Split_348_n804_AND2T_72_n96(net277_c1,net277);
INTERCONNECT Split_356_n812_OR2T_102_n126(net278_c1,net278);
INTERCONNECT Split_364_n820_DFFT_162__FBL_n618(net279_c1,net279);
INTERCONNECT Split_349_n805_DFFT_167__FBL_n623(net280_c1,net280);
INTERCONNECT Split_357_n813_OR2T_127_n151(net281_c1,net281);
INTERCONNECT Split_365_n821_Split_366_n822(net282_c1,net282);
INTERCONNECT Split_358_n814_OR2T_115_n139(net283_c1,net283);
INTERCONNECT Split_366_n822_AND2T_61_n85(net284_c1,net284);
INTERCONNECT Split_374_n830_XOR2T_45_n69(net285_c1,net285);
INTERCONNECT Split_350_n806_DFFT_159__FBL_n615(net286_c1,net286);
INTERCONNECT Split_359_n815_OR2T_115_n139(net287_c1,net287);
INTERCONNECT Split_367_n823_DFFT_187__FPB_n643(net288_c1,net288);
INTERCONNECT Split_375_n831_Split_376_n832(net289_c1,net289);
INTERCONNECT Split_351_n807_OR2T_93_n117(net290_c1,net290);
INTERCONNECT Split_368_n824_Split_369_n825(net291_c1,net291);
INTERCONNECT Split_376_n832_AND2T_26_n50(net292_c1,net292);
INTERCONNECT Split_384_n840_Split_385_n841(net293_c1,net293);
INTERCONNECT Split_352_n808_Split_353_n809(net294_c1,net294);
INTERCONNECT Split_360_n816_Split_361_n817(net295_c1,net295);
INTERCONNECT Split_369_n825_AND2T_16_n40(net296_c1,net296);
INTERCONNECT Split_377_n833_AND2T_39_n63(net297_c1,net297);
INTERCONNECT Split_385_n841_AND2T_51_n75(net298_c1,net298);
INTERCONNECT Split_353_n809_DFFT_160__FBL_n616(net299_c1,net299);
INTERCONNECT Split_361_n817_DFFT_161__FBL_n617(net300_c1,net300);
INTERCONNECT Split_378_n834_Split_379_n835(net301_c1,net301);
INTERCONNECT Split_386_n842_OR2T_58_n82(net302_c1,net302);
INTERCONNECT Split_394_n850_AND2T_18_n42(net303_c1,net303);
INTERCONNECT Split_362_n818_DFFT_169__FBL_n625(net304_c1,net304);
INTERCONNECT Split_370_n826_AND2T_68_n92(net305_c1,net305);
INTERCONNECT Split_314_n770_Split_315_n771(net306_c1,net306);
INTERCONNECT Split_379_n835_AND2T_29_n53(net307_c1,net307);
INTERCONNECT Split_387_n843_Split_388_n844(net308_c1,net308);
INTERCONNECT Split_395_n851_AND2T_85_n109(net309_c1,net309);
INTERCONNECT Split_363_n819_DFFT_170__FBL_n626(net310_c1,net310);
INTERCONNECT Split_371_n827_AND2T_143_n179(net311_c1,net311);
INTERCONNECT Split_307_n763_Split_308_n764(net312_c1,net312);
INTERCONNECT Split_315_n771_AND2T_15_n39(net313_c1,net313);
INTERCONNECT Split_388_n844_AND2T_85_n109(net314_c1,net314);
INTERCONNECT Split_396_n852_Split_397_n853(net315_c1,net315);
INTERCONNECT Split_372_n828_Split_373_n829(net316_c1,net316);
INTERCONNECT Split_380_n836_OR2T_42_n66(net317_c1,net317);
INTERCONNECT Split_308_n764_NOTT_147_n183(net318_c1,net318);
INTERCONNECT Split_316_n772_AND2T_141_n177(net319_c1,net319);
INTERCONNECT Split_324_n780_AND2T_87_n111(net320_c1,net320);
INTERCONNECT Split_404_n860_DFFT_257__FPB_n713(net321_c1,net321);
INTERCONNECT Split_389_n845_DFFT_230__FPB_n686(net322_c1,net322);
INTERCONNECT Split_397_n853_AND2T_21_n45(net323_c1,net323);
INTERCONNECT Split_373_n829_AND2T_22_n46(net324_c1,net324);
INTERCONNECT Split_381_n837_Split_382_n838(net325_c1,net325);
INTERCONNECT Split_309_n765_DFFT_152__FPB_n206(net326_c1,net326);
INTERCONNECT Split_317_n773_OR2T_23_n47(net327_c1,net327);
INTERCONNECT Split_325_n781_Split_326_n782(net328_c1,net328);
INTERCONNECT Split_405_n861_Split_406_n862(net329_c1,net329);
INTERCONNECT Split_398_n854_AND2T_90_n114(net330_c1,net330);
INTERCONNECT Split_382_n838_NOTT_41_n65(net331_c1,net331);
INTERCONNECT Split_390_n846_Split_391_n847(net332_c1,net332);
INTERCONNECT Split_318_n774_Split_319_n775(net333_c1,net333);
INTERCONNECT Split_326_n782_AND2T_26_n50(net334_c1,net334);
INTERCONNECT Split_334_n790_AND2T_133_n157(net335_c1,net335);
INTERCONNECT Split_406_n862_NOTT_8_n32(net336_c1,net336);
INTERCONNECT Split_414_n870_XOR2T_36_n60(net337_c1,net337);
INTERCONNECT Split_310_n766_NOTT_138_n162(net338_c1,net338);
INTERCONNECT Split_399_n855_Split_400_n856(net339_c1,net339);
INTERCONNECT Split_383_n839_DFFT_186__FPB_n642(net340_c1,net340);
INTERCONNECT Split_391_n847_AND2T_21_n45(net341_c1,net341);
INTERCONNECT Split_319_n775_AND2T_22_n46(net342_c1,net342);
INTERCONNECT Split_327_n783_AND2T_52_n76(net343_c1,net343);
INTERCONNECT Split_335_n791_OR2T_34_n58(net344_c1,net344);
INTERCONNECT Split_407_n863_NOTT_97_n121(net345_c1,net345);
INTERCONNECT Split_415_n871_NOTT_149_n197(net346_c1,net346);
INTERCONNECT Split_311_n767_Split_312_n768(net347_c1,net347);
INTERCONNECT Split_392_n848_AND2T_67_n91(net348_c1,net348);
INTERCONNECT Split_328_n784_OR2T_30_n54(net349_c1,net349);
INTERCONNECT Split_336_n792_NOTT_40_n64(net350_c1,net350);
INTERCONNECT Split_408_n864_DFFT_203__FPB_n659(net351_c1,net351);
INTERCONNECT Split_416_n872_AND2T_140_n176(net352_c1,net352);
INTERCONNECT Split_424_n880_NOTT_14_n38(net353_c1,net353);
INTERCONNECT Split_312_n768_AND2T_9_n33(net354_c1,net354);
INTERCONNECT Split_320_n776_AND2T_66_n90(net355_c1,net355);
INTERCONNECT Split_400_n856_NOTT_50_n74(net356_c1,net356);
INTERCONNECT Split_393_n849_Split_394_n850(net357_c1,net357);
INTERCONNECT Split_329_n785_AND2T_113_n137(net358_c1,net358);
INTERCONNECT Split_337_n793_OR2T_42_n66(net359_c1,net359);
INTERCONNECT Split_409_n865_DFFT_195__FPB_n651(net360_c1,net360);
INTERCONNECT Split_417_n873_AND2T_140_n176(net361_c1,net361);
INTERCONNECT Split_425_n881_DFFT_179__FPB_n635(net362_c1,net362);
INTERCONNECT Split_313_n769_AND2T_11_n35(net363_c1,net363);
INTERCONNECT Split_321_n777_AND2T_106_n130(net364_c1,net364);
INTERCONNECT Split_401_n857_AND2T_90_n114(net365_c1,net365);
INTERCONNECT Split_338_n794_AND2T_46_n70(net366_c1,net366);
INTERCONNECT Split_418_n874_AND2T_146_n182(net367_c1,net367);
INTERCONNECT Split_426_n882_Split_427_n883(net368_c1,net368);
INTERCONNECT Split_322_n778_OR2T_23_n47(net369_c1,net369);
INTERCONNECT Split_330_n786_AND2T_71_n95(net370_c1,net370);
INTERCONNECT Split_402_n858_Split_403_n859(net371_c1,net371);
INTERCONNECT Split_410_n866_DFFT_241__FPB_n697(net372_c1,net372);
INTERCONNECT Split_339_n795_Split_340_n796(net373_c1,net373);
INTERCONNECT Split_419_n875_AND2T_146_n182(net374_c1,net374);
INTERCONNECT Split_427_n883_AND2T_13_n37(net375_c1,net375);
INTERCONNECT Split_323_n779_OR2T_127_n151(net376_c1,net376);
INTERCONNECT Split_331_n787_DFFT_209__FPB_n665(net377_c1,net377);
INTERCONNECT Split_403_n859_AND2T_101_n125(net378_c1,net378);
INTERCONNECT Split_411_n867_AND2T_84_n108(net379_c1,net379);
INTERCONNECT Split_428_n884_DFFT_175__FPB_n631(net380_c1,net380);
INTERCONNECT Split_332_n788_OR2T_30_n54(net381_c1,net381);
INTERCONNECT Split_340_n796_OR2T_78_n102(net382_c1,net382);
INTERCONNECT Split_412_n868_DFFT_244__FPB_n700(net383_c1,net383);
INTERCONNECT Split_420_n876_Split_421_n877(net384_c1,net384);
INTERCONNECT Split_429_n885_Split_430_n886(net385_c1,net385);
INTERCONNECT Split_333_n789_OR2T_34_n58(net386_c1,net386);
INTERCONNECT Split_341_n797_OR2T_119_n143(net387_c1,net387);
INTERCONNECT Split_413_n869_XOR2T_36_n60(net388_c1,net388);
INTERCONNECT Split_421_n877_AND2T_13_n37(net389_c1,net389);
INTERCONNECT Split_342_n798_AND2T_123_n147(net390_c1,net390);
INTERCONNECT Split_422_n878_DFFT_173__FPB_n629(net391_c1,net391);
INTERCONNECT Split_430_n886_NOTT_17_n41(net392_c1,net392);
INTERCONNECT Split_343_n799_DFFT_212__FPB_n668(net393_c1,net393);
INTERCONNECT Split_423_n879_Split_424_n880(net394_c1,net394);
INTERCONNECT Split_431_n887_DFFT_177__FPB_n633(net395_c1,net395);
INTERCONNECT DFFT_156__PIPL_n210_DFFT_286__FPB_n742(net396_c1,net396);
INTERCONNECT DFFT_157__PIPL_n211_DFFT_293__FPB_n749(net397_c1,net397);
INTERCONNECT DFFT_158__PIPL_n212_DFFT_300__FPB_n756(net398_c1,net398);
INTERCONNECT DFFT_155__PIPL_n209_Split_HOLD_944(net399_c1,net399);
INTERCONNECT DFFT_164__FBL_n620_Split_417_n873(net400_c1,net400);
INTERCONNECT DFFT_165__FBL_n621_Split_418_n874(net401_c1,net401);
INTERCONNECT DFFT_166__FBL_n622_Split_419_n875(net402_c1,net402);
INTERCONNECT DFFT_167__FBL_n623_Split_420_n876(net403_c1,net403);
INTERCONNECT DFFT_159__FBL_n615_Split_408_n864(net404_c1,net404);
INTERCONNECT DFFT_160__FBL_n616_Split_410_n866(net405_c1,net405);
INTERCONNECT DFFT_168__FBL_n624_NOTT_151_n199(net406_c1,net406);
INTERCONNECT DFFT_161__FBL_n617_Split_412_n868(net407_c1,net407);
INTERCONNECT DFFT_169__FBL_n625_Split_HOLD_943(net408_c1,net408);
INTERCONNECT DFFT_170__FBL_n626_Split_423_n879(net409_c1,net409);
INTERCONNECT DFFT_162__FBL_n618_Split_414_n870(net410_c1,net410);
INTERCONNECT DFFT_171__FBL_n627_Split_426_n882(net411_c1,net411);
INTERCONNECT DFFT_163__FBL_n619_Split_415_n871(net412_c1,net412);
INTERCONNECT DFFT_172__FBL_n628_Split_429_n885(net413_c1,net413);
INTERCONNECT DFFT_152__FPB_n206_Split_399_n855(net414_c1,net414);
INTERCONNECT DFFT_153__FPB_n207_Split_402_n858(net415_c1,net415);
INTERCONNECT DFFT_154__FPB_n208_Split_405_n861(net416_c1,net416);
INTERCONNECT DFFT_244__FPB_n700_AND2T_105_n129(net417_c1,net417);
INTERCONNECT DFFT_245__FPB_n701_AND2T_106_n130(net418_c1,net418);
INTERCONNECT DFFT_254__FPB_n710_DFFT_255__FPB_n711(net419_c1,net419);
INTERCONNECT DFFT_246__FPB_n702_OR2T_108_n132(net420_c1,net420);
INTERCONNECT DFFT_174__FPB_n630_AND2T_9_n33(net421_c1,net421);
INTERCONNECT DFFT_255__FPB_n711_DFFT_256__FPB_n712(net422_c1,net422);
INTERCONNECT DFFT_175__FPB_n631_DFFT_176__FPB_n632(net423_c1,net423);
INTERCONNECT DFFT_247__FPB_n703_AND2T_109_n133(net424_c1,net424);
INTERCONNECT DFFT_264__FPB_n720_AND2T_132_n156(net425_c1,net425);
INTERCONNECT DFFT_256__FPB_n712_AND2T_121_n145(net426_c1,net426);
INTERCONNECT DFFT_248__FPB_n704_OR2T_112_n136(net427_c1,net427);
INTERCONNECT DFFT_184__FPB_n640_AND2T_25_n49(net428_c1,net428);
INTERCONNECT DFFT_176__FPB_n632_AND2T_10_n34(net429_c1,net429);
INTERCONNECT DFFT_265__FPB_n721_DFFT_266__FPB_n722(net430_c1,net430);
INTERCONNECT DFFT_257__FPB_n713_DFFT_258__FPB_n714(net431_c1,net431);
INTERCONNECT DFFT_177__FPB_n633_DFFT_178__FPB_n634(net432_c1,net432);
INTERCONNECT DFFT_249__FPB_n705_OR2T_119_n143(net433_c1,net433);
INTERCONNECT DFFT_185__FPB_n641_AND2T_27_n51(net434_c1,net434);
INTERCONNECT DFFT_274__FPB_n730_DFFT_275__FPB_n731(net435_c1,net435);
INTERCONNECT DFFT_250__FPB_n706_DFFT_251__FPB_n707(net436_c1,net436);
INTERCONNECT DFFT_266__FPB_n722_AND2T_133_n157(net437_c1,net437);
INTERCONNECT DFFT_258__FPB_n714_AND2T_122_n146(net438_c1,net438);
INTERCONNECT DFFT_194__FPB_n650_AND2T_48_n72(net439_c1,net439);
INTERCONNECT DFFT_186__FPB_n642_AND2T_29_n53(net440_c1,net440);
INTERCONNECT DFFT_178__FPB_n634_AND2T_11_n35(net441_c1,net441);
INTERCONNECT DFFT_259__FPB_n715_DFFT_260__FPB_n716(net442_c1,net442);
INTERCONNECT DFFT_251__FPB_n707_DFFT_252__FPB_n708(net443_c1,net443);
INTERCONNECT DFFT_179__FPB_n635_DFFT_180__FPB_n636(net444_c1,net444);
INTERCONNECT DFFT_275__FPB_n731_AND2T_139_n163(net445_c1,net445);
INTERCONNECT DFFT_267__FPB_n723_OR2T_137_n161(net446_c1,net446);
INTERCONNECT DFFT_195__FPB_n651_AND2T_51_n75(net447_c1,net447);
INTERCONNECT DFFT_187__FPB_n643_AND2T_32_n56(net448_c1,net448);
INTERCONNECT DFFT_284__FPB_n740_DFFT_285_state_obs0(net449_c1,net449);
INTERCONNECT DFFT_268__FPB_n724_DFFT_269__FPB_n725(net450_c1,net450);
INTERCONNECT DFFT_252__FPB_n708_DFFT_253__FPB_n709(net451_c1,net451);
INTERCONNECT DFFT_276__FPB_n732_AND2T_141_n177(net452_c1,net452);
INTERCONNECT DFFT_260__FPB_n716_AND2T_123_n147(net453_c1,net453);
INTERCONNECT DFFT_204__FPB_n660_OR2T_60_n84(net454_c1,net454);
INTERCONNECT DFFT_196__FPB_n652_AND2T_52_n76(net455_c1,net455);
INTERCONNECT DFFT_188__FPB_n644_AND2T_35_n59(net456_c1,net456);
INTERCONNECT DFFT_180__FPB_n636_AND2T_12_n36(net457_c1,net457);
INTERCONNECT DFFT_269__FPB_n725_DFFT_270__FPB_n726(net458_c1,net458);
INTERCONNECT DFFT_253__FPB_n709_DFFT_254__FPB_n710(net459_c1,net459);
INTERCONNECT DFFT_173__FPB_n629_DFFT_174__FPB_n630(net460_c1,net460);
INTERCONNECT DFFT_277__FPB_n733_AND2T_144_n180(net461_c1,net461);
INTERCONNECT DFFT_261__FPB_n717_AND2T_124_n148(net462_c1,net462);
INTERCONNECT DFFT_205__FPB_n661_OR2T_62_n86(net463_c1,net463);
INTERCONNECT DFFT_197__FPB_n653_AND2T_53_n77(net464_c1,net464);
INTERCONNECT DFFT_189__FPB_n645_OR2T_37_n61(net465_c1,net465);
INTERCONNECT DFFT_181__FPB_n637_AND2T_15_n39(net466_c1,net466);
INTERCONNECT DFFT_294__FPB_n750_DFFT_295__FPB_n751(net467_c1,net467);
INTERCONNECT DFFT_286__FPB_n742_DFFT_287__FPB_n743(net468_c1,net468);
INTERCONNECT DFFT_270__FPB_n726_DFFT_271__FPB_n727(net469_c1,net469);
INTERCONNECT DFFT_206__FPB_n662_DFFT_207__FPB_n663(net470_c1,net470);
INTERCONNECT DFFT_198__FPB_n654_DFFT_199__FPB_n655(net471_c1,net471);
INTERCONNECT DFFT_278__FPB_n734_AND2T_145_n181(net472_c1,net472);
INTERCONNECT DFFT_262__FPB_n718_OR2T_126_n150(net473_c1,net473);
INTERCONNECT DFFT_214__FPB_n670_OR2T_77_n101(net474_c1,net474);
INTERCONNECT DFFT_190__FPB_n646_AND2T_43_n67(net475_c1,net475);
INTERCONNECT DFFT_182__FPB_n638_AND2T_16_n40(net476_c1,net476);
INTERCONNECT DFFT_295__FPB_n751_DFFT_296__FPB_n752(net477_c1,net477);
INTERCONNECT DFFT_287__FPB_n743_DFFT_288__FPB_n744(net478_c1,net478);
INTERCONNECT DFFT_279__FPB_n735_DFFT_280__FPB_n736(net479_c1,net479);
INTERCONNECT DFFT_271__FPB_n727_DFFT_272__FPB_n728(net480_c1,net480);
INTERCONNECT DFFT_215__FPB_n671_DFFT_216__FPB_n672(net481_c1,net481);
INTERCONNECT DFFT_207__FPB_n663_DFFT_208__FPB_n664(net482_c1,net482);
INTERCONNECT DFFT_191__FPB_n647_DFFT_192__FPB_n648(net483_c1,net483);
INTERCONNECT DFFT_263__FPB_n719_AND2T_128_n152(net484_c1,net484);
INTERCONNECT DFFT_199__FPB_n655_AND2T_54_n78(net485_c1,net485);
INTERCONNECT DFFT_183__FPB_n639_AND2T_24_n48(net486_c1,net486);
INTERCONNECT DFFT_304__FPB_n760_DFFT_305__FPB_n761(net487_c1,net487);
INTERCONNECT DFFT_296__FPB_n752_DFFT_297__FPB_n753(net488_c1,net488);
INTERCONNECT DFFT_288__FPB_n744_DFFT_289__FPB_n745(net489_c1,net489);
INTERCONNECT DFFT_280__FPB_n736_DFFT_281__FPB_n737(net490_c1,net490);
INTERCONNECT DFFT_272__FPB_n728_DFFT_273__FPB_n729(net491_c1,net491);
INTERCONNECT DFFT_224__FPB_n680_DFFT_225__FPB_n681(net492_c1,net492);
INTERCONNECT DFFT_216__FPB_n672_DFFT_217__FPB_n673(net493_c1,net493);
INTERCONNECT DFFT_208__FPB_n664_AND2T_63_n87(net494_c1,net494);
INTERCONNECT DFFT_200__FPB_n656_XOR2T_55_n79(net495_c1,net495);
INTERCONNECT DFFT_192__FPB_n648_AND2T_44_n68(net496_c1,net496);
INTERCONNECT DFFT_305__FPB_n761_DFFT_306_state_obs3(net497_c1,net497);
INTERCONNECT DFFT_297__FPB_n753_DFFT_298__FPB_n754(net498_c1,net498);
INTERCONNECT DFFT_289__FPB_n745_DFFT_290__FPB_n746(net499_c1,net499);
INTERCONNECT DFFT_281__FPB_n737_DFFT_282__FPB_n738(net500_c1,net500);
INTERCONNECT DFFT_273__FPB_n729_DFFT_274__FPB_n730(net501_c1,net501);
INTERCONNECT DFFT_225__FPB_n681_DFFT_226__FPB_n682(net502_c1,net502);
INTERCONNECT DFFT_217__FPB_n673_DFFT_218__FPB_n674(net503_c1,net503);
INTERCONNECT DFFT_209__FPB_n665_AND2T_64_n88(net504_c1,net504);
INTERCONNECT DFFT_201__FPB_n657_AND2T_56_n80(net505_c1,net505);
INTERCONNECT DFFT_193__FPB_n649_Split_HOLD_945(net506_c1,net506);
INTERCONNECT DFFT_298__FPB_n754_DFFT_299_state_obs2(net507_c1,net507);
INTERCONNECT DFFT_290__FPB_n746_DFFT_291__FPB_n747(net508_c1,net508);
INTERCONNECT DFFT_282__FPB_n738_DFFT_283__FPB_n739(net509_c1,net509);
INTERCONNECT DFFT_234__FPB_n690_DFFT_235__FPB_n691(net510_c1,net510);
INTERCONNECT DFFT_218__FPB_n674_DFFT_219__FPB_n675(net511_c1,net511);
INTERCONNECT DFFT_210__FPB_n666_DFFT_211__FPB_n667(net512_c1,net512);
INTERCONNECT DFFT_226__FPB_n682_AND2T_81_n105(net513_c1,net513);
INTERCONNECT DFFT_202__FPB_n658_AND2T_57_n81(net514_c1,net514);
INTERCONNECT DFFT_291__FPB_n747_DFFT_292_state_obs1(net515_c1,net515);
INTERCONNECT DFFT_283__FPB_n739_DFFT_284__FPB_n740(net516_c1,net516);
INTERCONNECT DFFT_235__FPB_n691_DFFT_236__FPB_n692(net517_c1,net517);
INTERCONNECT DFFT_227__FPB_n683_DFFT_228__FPB_n684(net518_c1,net518);
INTERCONNECT DFFT_219__FPB_n675_DFFT_220__FPB_n676(net519_c1,net519);
INTERCONNECT DFFT_211__FPB_n667_AND2T_72_n96(net520_c1,net520);
INTERCONNECT DFFT_203__FPB_n659_OR2T_58_n82(net521_c1,net521);
INTERCONNECT DFFT_300__FPB_n756_DFFT_301__FPB_n757(net522_c1,net522);
INTERCONNECT DFFT_236__FPB_n692_DFFT_237__FPB_n693(net523_c1,net523);
INTERCONNECT DFFT_220__FPB_n676_DFFT_221__FPB_n677(net524_c1,net524);
INTERCONNECT DFFT_228__FPB_n684_OR2T_89_n113(net525_c1,net525);
INTERCONNECT DFFT_212__FPB_n668_AND2T_73_n97(net526_c1,net526);
INTERCONNECT DFFT_301__FPB_n757_DFFT_302__FPB_n758(net527_c1,net527);
INTERCONNECT DFFT_293__FPB_n749_DFFT_294__FPB_n750(net528_c1,net528);
INTERCONNECT DFFT_237__FPB_n693_DFFT_238__FPB_n694(net529_c1,net529);
INTERCONNECT DFFT_229__FPB_n685_AND2T_91_n115(net530_c1,net530);
INTERCONNECT DFFT_221__FPB_n677_AND2T_80_n104(net531_c1,net531);
INTERCONNECT DFFT_213__FPB_n669_OR2T_76_n100(net532_c1,net532);
INTERCONNECT DFFT_302__FPB_n758_DFFT_303__FPB_n759(net533_c1,net533);
INTERCONNECT DFFT_238__FPB_n694_DFFT_239__FPB_n695(net534_c1,net534);
INTERCONNECT DFFT_230__FPB_n686_DFFT_231__FPB_n687(net535_c1,net535);
INTERCONNECT DFFT_222__FPB_n678_DFFT_223__FPB_n679(net536_c1,net536);
INTERCONNECT DFFT_303__FPB_n759_DFFT_304__FPB_n760(net537_c1,net537);
INTERCONNECT DFFT_223__FPB_n679_DFFT_224__FPB_n680(net538_c1,net538);
INTERCONNECT DFFT_239__FPB_n695_AND2T_98_n122(net539_c1,net539);
INTERCONNECT DFFT_231__FPB_n687_AND2T_92_n116(net540_c1,net540);
INTERCONNECT DFFT_240__FPB_n696_AND2T_99_n123(net541_c1,net541);
INTERCONNECT DFFT_232__FPB_n688_OR2T_95_n119(net542_c1,net542);
INTERCONNECT DFFT_233__FPB_n689_DFFT_234__FPB_n690(net543_c1,net543);
INTERCONNECT DFFT_241__FPB_n697_AND2T_101_n125(net544_c1,net544);
INTERCONNECT DFFT_242__FPB_n698_DFFT_243__FPB_n699(net545_c1,net545);
INTERCONNECT DFFT_243__FPB_n699_AND2T_104_n128(net546_c1,net546);
INTERCONNECT DFFT_285_state_obs0_state_obs0_Pad(net547_c1,state_obs0_Pad);
INTERCONNECT DFFT_292_state_obs1_state_obs1_Pad(net548_c1,state_obs1_Pad);
INTERCONNECT DFFT_299_state_obs2_state_obs2_Pad(net549_c1,state_obs2_Pad);
INTERCONNECT DFFT_306_state_obs3_state_obs3_Pad(net550_c1,state_obs3_Pad);
INTERCONNECT SplitCLK_0_810_SplitCLK_0_448(net551_c1,net551);
INTERCONNECT SplitCLK_0_810_SplitCLK_2_596(net552_c1,net552);
INTERCONNECT SplitCLK_2_809_DFFT_198__FPB_n654(net553_c1,net553);
INTERCONNECT SplitCLK_2_808_DFFT_278__FPB_n734(net554_c1,net554);
INTERCONNECT SplitCLK_4_807_DFFT_286__FPB_n742(net555_c1,net555);
INTERCONNECT SplitCLK_4_806_DFFT_294__FPB_n750(net556_c1,net556);
INTERCONNECT SplitCLK_2_805_DFFT_293__FPB_n749(net557_c1,net557);
INTERCONNECT SplitCLK_4_804_DFFT_197__FPB_n653(net558_c1,net558);
INTERCONNECT SplitCLK_2_803_DFFT_269__FPB_n725(net559_c1,net559);
INTERCONNECT SplitCLK_4_802_DFFT_277__FPB_n733(net560_c1,net560);
INTERCONNECT SplitCLK_2_801_NOTT_97_n121(net561_c1,net561);
INTERCONNECT SplitCLK_2_800_NOTT_79_n103(net562_c1,net562);
INTERCONNECT SplitCLK_4_799_DFFT_188__FPB_n644(net563_c1,net563);
INTERCONNECT SplitCLK_2_798_DFFT_196__FPB_n652(net564_c1,net564);
INTERCONNECT SplitCLK_4_797_DFFT_268__FPB_n724(net565_c1,net565);
INTERCONNECT SplitCLK_4_796_DFFT_276__FPB_n732(net566_c1,net566);
INTERCONNECT SplitCLK_4_795_NOTT_82_n106(net567_c1,net567);
INTERCONNECT SplitCLK_2_794_DFFT_179__FPB_n635(net568_c1,net568);
INTERCONNECT SplitCLK_2_793_DFFT_187__FPB_n643(net569_c1,net569);
INTERCONNECT SplitCLK_4_792_DFFT_195__FPB_n651(net570_c1,net570);
INTERCONNECT SplitCLK_4_791_DFFT_259__FPB_n715(net571_c1,net571);
INTERCONNECT SplitCLK_2_790_DFFT_267__FPB_n723(net572_c1,net572);
INTERCONNECT SplitCLK_2_789_DFFT_275__FPB_n731(net573_c1,net573);
INTERCONNECT SplitCLK_2_788_DFFT_282__FPB_n738(net574_c1,net574);
INTERCONNECT SplitCLK_2_787_DFFT_178__FPB_n634(net575_c1,net575);
INTERCONNECT SplitCLK_4_786_DFFT_186__FPB_n642(net576_c1,net576);
INTERCONNECT SplitCLK_4_785_DFFT_194__FPB_n650(net577_c1,net577);
INTERCONNECT SplitCLK_4_784_DFFT_274__FPB_n730(net578_c1,net578);
INTERCONNECT SplitCLK_4_783_DFFT_193__FPB_n649(net579_c1,net579);
INTERCONNECT SplitCLK_2_782_DFFT_273__FPB_n729(net580_c1,net580);
INTERCONNECT SplitCLK_4_781_DFFT_281__FPB_n737(net581_c1,net581);
INTERCONNECT SplitCLK_4_780_DFFT_177__FPB_n633(net582_c1,net582);
INTERCONNECT SplitCLK_4_779_DFFT_185__FPB_n641(net583_c1,net583);
INTERCONNECT SplitCLK_4_778_DFFT_257__FPB_n713(net584_c1,net584);
INTERCONNECT SplitCLK_2_777_DFFT_192__FPB_n648(net585_c1,net585);
INTERCONNECT SplitCLK_4_776_DFFT_272__FPB_n728(net586_c1,net586);
INTERCONNECT SplitCLK_2_775_DFFT_280__FPB_n736(net587_c1,net587);
INTERCONNECT SplitCLK_2_774_DFFT_176__FPB_n632(net588_c1,net588);
INTERCONNECT SplitCLK_4_773_DFFT_248__FPB_n704(net589_c1,net589);
INTERCONNECT SplitCLK_4_772_DFFT_256__FPB_n712(net590_c1,net590);
INTERCONNECT SplitCLK_4_771_NOTT_148_n184(net591_c1,net591);
INTERCONNECT SplitCLK_4_770_NOTT_147_n183(net592_c1,net592);
INTERCONNECT SplitCLK_2_769_NOTT_138_n162(net593_c1,net593);
INTERCONNECT SplitCLK_4_768_NOTT_151_n199(net594_c1,net594);
INTERCONNECT SplitCLK_2_767_NOTT_142_n178(net595_c1,net595);
INTERCONNECT SplitCLK_4_766_DFFT_168__FBL_n624(net596_c1,net596);
INTERCONNECT SplitCLK_4_765_DFFT_239__FPB_n695(net597_c1,net597);
INTERCONNECT SplitCLK_2_764_DFFT_183__FPB_n639(net598_c1,net598);
INTERCONNECT SplitCLK_4_763_DFFT_191__FPB_n647(net599_c1,net599);
INTERCONNECT SplitCLK_2_762_DFFT_263__FPB_n719(net600_c1,net600);
INTERCONNECT SplitCLK_2_761_DFFT_271__FPB_n727(net601_c1,net601);
INTERCONNECT SplitCLK_2_760_DFFT_247__FPB_n703(net602_c1,net602);
INTERCONNECT SplitCLK_4_759_DFFT_255__FPB_n711(net603_c1,net603);
INTERCONNECT SplitCLK_4_758_DFFT_159__FBL_n615(net604_c1,net604);
INTERCONNECT SplitCLK_2_757_DFFT_238__FPB_n694(net605_c1,net605);
INTERCONNECT SplitCLK_4_756_DFFT_182__FPB_n638(net606_c1,net606);
INTERCONNECT SplitCLK_4_755_DFFT_270__FPB_n726(net607_c1,net607);
INTERCONNECT SplitCLK_2_754_DFFT_246__FPB_n702(net608_c1,net608);
INTERCONNECT SplitCLK_4_753_DFFT_166__FBL_n622(net609_c1,net609);
INTERCONNECT SplitCLK_2_752_DFFT_229__FPB_n685(net610_c1,net610);
INTERCONNECT SplitCLK_4_751_DFFT_237__FPB_n693(net611_c1,net611);
INTERCONNECT SplitCLK_4_750_DFFT_173__FPB_n629(net612_c1,net612);
INTERCONNECT SplitCLK_2_749_DFFT_181__FPB_n637(net613_c1,net613);
INTERCONNECT SplitCLK_4_748_DFFT_165__FBL_n621(net614_c1,net614);
INTERCONNECT SplitCLK_4_747_DFFT_236__FPB_n692(net615_c1,net615);
INTERCONNECT SplitCLK_4_746_DFFT_180__FPB_n636(net616_c1,net616);
INTERCONNECT SplitCLK_2_745_DFFT_252__FPB_n708(net617_c1,net617);
INTERCONNECT SplitCLK_4_744_DFFT_260__FPB_n716(net618_c1,net618);
INTERCONNECT SplitCLK_4_743_DFFT_244__FPB_n700(net619_c1,net619);
INTERCONNECT SplitCLK_4_742_DFFT_164__FBL_n620(net620_c1,net620);
INTERCONNECT SplitCLK_2_741_DFFT_219__FPB_n675(net621_c1,net621);
INTERCONNECT SplitCLK_4_740_DFFT_251__FPB_n707(net622_c1,net622);
INTERCONNECT SplitCLK_2_739_DFFT_163__FBL_n619(net623_c1,net623);
INTERCONNECT SplitCLK_2_738_DFFT_242__FPB_n698(net624_c1,net624);
INTERCONNECT SplitCLK_4_737_DFFT_218__FPB_n674(net625_c1,net625);
INTERCONNECT SplitCLK_2_736_DFFT_226__FPB_n682(net626_c1,net626);
INTERCONNECT SplitCLK_2_735_DFFT_250__FPB_n706(net627_c1,net627);
INTERCONNECT SplitCLK_4_734_DFFT_154__FPB_n208(net628_c1,net628);
INTERCONNECT SplitCLK_4_733_DFFT_162__FBL_n618(net629_c1,net629);
INTERCONNECT SplitCLK_4_732_DFFT_170__FBL_n626(net630_c1,net630);
INTERCONNECT SplitCLK_2_731_DFFT_233__FPB_n689(net631_c1,net631);
INTERCONNECT SplitCLK_4_730_DFFT_209__FPB_n665(net632_c1,net632);
INTERCONNECT SplitCLK_4_729_DFFT_217__FPB_n673(net633_c1,net633);
INTERCONNECT SplitCLK_4_728_DFFT_225__FPB_n681(net634_c1,net634);
INTERCONNECT SplitCLK_2_727_DFFT_305__FPB_n761(net635_c1,net635);
INTERCONNECT SplitCLK_2_726_OR2T_89_n113(net636_c1,net636);
INTERCONNECT SplitCLK_4_725_OR2T_96_n120(net637_c1,net637);
INTERCONNECT SplitCLK_4_724_DFFT_232__FPB_n688(net638_c1,net638);
INTERCONNECT SplitCLK_4_723_OR2T_95_n119(net639_c1,net639);
INTERCONNECT SplitCLK_4_722_DFFT_208__FPB_n664(net640_c1,net640);
INTERCONNECT SplitCLK_2_721_DFFT_216__FPB_n672(net641_c1,net641);
INTERCONNECT SplitCLK_2_720_DFFT_224__FPB_n680(net642_c1,net642);
INTERCONNECT SplitCLK_4_719_DFFT_304__FPB_n760(net643_c1,net643);
INTERCONNECT SplitCLK_4_718_OR2T_94_n118(net644_c1,net644);
INTERCONNECT SplitCLK_2_717_DFFT_152__FPB_n206(net645_c1,net645);
INTERCONNECT SplitCLK_2_716_OR2T_78_n102(net646_c1,net646);
INTERCONNECT SplitCLK_4_715_OR2T_93_n117(net647_c1,net647);
INTERCONNECT SplitCLK_4_714_DFFT_158__PIPL_n212(net648_c1,net648);
INTERCONNECT SplitCLK_4_713_OR2T_76_n100(net649_c1,net649);
INTERCONNECT SplitCLK_2_712_DFFT_231__FPB_n687(net650_c1,net650);
INTERCONNECT SplitCLK_2_711_DFFT_207__FPB_n663(net651_c1,net651);
INTERCONNECT SplitCLK_4_710_DFFT_215__FPB_n671(net652_c1,net652);
INTERCONNECT SplitCLK_4_709_DFFT_222__FPB_n678(net653_c1,net653);
INTERCONNECT SplitCLK_4_708_DFFT_230__FPB_n686(net654_c1,net654);
INTERCONNECT SplitCLK_4_707_DFFT_206__FPB_n662(net655_c1,net655);
INTERCONNECT SplitCLK_2_706_DFFT_214__FPB_n670(net656_c1,net656);
INTERCONNECT SplitCLK_4_705_DFFT_213__FPB_n669(net657_c1,net657);
INTERCONNECT SplitCLK_4_704_DFFT_212__FPB_n668(net658_c1,net658);
INTERCONNECT SplitCLK_2_703_DFFT_204__FPB_n660(net659_c1,net659);
INTERCONNECT SplitCLK_2_702_DFFT_156__PIPL_n210(net660_c1,net660);
INTERCONNECT SplitCLK_4_701_DFFT_203__FPB_n659(net661_c1,net661);
INTERCONNECT SplitCLK_2_700_DFFT_202__FPB_n658(net662_c1,net662);
INTERCONNECT SplitCLK_4_699_DFFT_210__FPB_n666(net663_c1,net663);
INTERCONNECT SplitCLK_4_698_DFFT_155__PIPL_n209(net664_c1,net664);
INTERCONNECT SplitCLK_2_697_DFFT_201__FPB_n657(net665_c1,net665);
INTERCONNECT SplitCLK_4_696_DFFT_200__FPB_n656(net666_c1,net666);
INTERCONNECT SplitCLK_2_695_AND2T_99_n123(net667_c1,net667);
INTERCONNECT SplitCLK_2_694_AND2T_87_n111(net668_c1,net668);
INTERCONNECT SplitCLK_2_693_AND2T_85_n109(net669_c1,net669);
INTERCONNECT SplitCLK_4_692_AND2T_84_n108(net670_c1,net670);
INTERCONNECT SplitCLK_4_691_AND2T_92_n116(net671_c1,net671);
INTERCONNECT SplitCLK_4_690_AND2T_83_n107(net672_c1,net672);
INTERCONNECT SplitCLK_2_689_AND2T_91_n115(net673_c1,net673);
INTERCONNECT SplitCLK_2_688_AND2T_81_n105(net674_c1,net674);
INTERCONNECT SplitCLK_2_687_AND2T_80_n104(net675_c1,net675);
INTERCONNECT SplitCLK_2_686_DFFT_299_state_obs2(net676_c1,net676);
INTERCONNECT SplitCLK_2_685_OR2T_137_n161(net677_c1,net677);
INTERCONNECT SplitCLK_4_684_OR2T_136_n160(net678_c1,net678);
INTERCONNECT SplitCLK_2_683_OR2T_135_n159(net679_c1,net679);
INTERCONNECT SplitCLK_4_682_OR2T_119_n143(net680_c1,net680);
INTERCONNECT SplitCLK_2_681_OR2T_127_n151(net681_c1,net681);
INTERCONNECT SplitCLK_2_680_OR2T_118_n142(net682_c1,net682);
INTERCONNECT SplitCLK_4_679_OR2T_125_n149(net683_c1,net683);
INTERCONNECT SplitCLK_2_678_OR2T_117_n141(net684_c1,net684);
INTERCONNECT SplitCLK_2_677_OR2T_108_n132(net685_c1,net685);
INTERCONNECT SplitCLK_4_676_OR2T_112_n136(net686_c1,net686);
INTERCONNECT SplitCLK_4_675_OR2T_102_n126(net687_c1,net687);
INTERCONNECT SplitCLK_4_674_NOTT_49_n73(net688_c1,net688);
INTERCONNECT SplitCLK_4_673_NOTT_47_n71(net689_c1,net689);
INTERCONNECT SplitCLK_4_672_NOTT_19_n43(net690_c1,net690);
INTERCONNECT SplitCLK_2_671_NOTT_50_n74(net691_c1,net691);
INTERCONNECT SplitCLK_2_670_NOTT_41_n65(net692_c1,net692);
INTERCONNECT SplitCLK_4_669_NOTT_17_n41(net693_c1,net693);
INTERCONNECT SplitCLK_4_668_NOTT_40_n64(net694_c1,net694);
INTERCONNECT SplitCLK_2_667_NOTT_14_n38(net695_c1,net695);
INTERCONNECT SplitCLK_4_666_NOTT_20_n44(net696_c1,net696);
INTERCONNECT SplitCLK_2_665_DFFT_285_state_obs0(net697_c1,net697);
INTERCONNECT SplitCLK_2_664_OR2T_75_n99(net698_c1,net698);
INTERCONNECT SplitCLK_2_663_OR2T_59_n83(net699_c1,net699);
INTERCONNECT SplitCLK_2_662_OR2T_74_n98(net700_c1,net700);
INTERCONNECT SplitCLK_4_661_OR2T_58_n82(net701_c1,net701);
INTERCONNECT SplitCLK_2_660_OR2T_65_n89(net702_c1,net702);
INTERCONNECT SplitCLK_2_659_OR2T_62_n86(net703_c1,net703);
INTERCONNECT SplitCLK_2_658_OR2T_70_n94(net704_c1,net704);
INTERCONNECT SplitCLK_2_657_OR2T_38_n62(net705_c1,net705);
INTERCONNECT SplitCLK_4_656_OR2T_60_n84(net706_c1,net706);
INTERCONNECT SplitCLK_2_655_OR2T_34_n58(net707_c1,net707);
INTERCONNECT SplitCLK_4_654_OR2T_42_n66(net708_c1,net708);
INTERCONNECT SplitCLK_4_653_OR2T_31_n55(net709_c1,net709);
INTERCONNECT SplitCLK_4_652_AND2T_68_n92(net710_c1,net710);
INTERCONNECT SplitCLK_2_651_AND2T_67_n91(net711_c1,net711);
INTERCONNECT SplitCLK_4_650_AND2T_66_n90(net712_c1,net712);
INTERCONNECT SplitCLK_2_649_AND2T_57_n81(net713_c1,net713);
INTERCONNECT SplitCLK_2_648_AND2T_64_n88(net714_c1,net714);
INTERCONNECT SplitCLK_4_647_AND2T_72_n96(net715_c1,net715);
INTERCONNECT SplitCLK_2_646_AND2T_48_n72(net716_c1,net716);
INTERCONNECT SplitCLK_2_645_AND2T_63_n87(net717_c1,net717);
INTERCONNECT SplitCLK_2_644_AND2T_71_n95(net718_c1,net718);
INTERCONNECT SplitCLK_4_643_AND2T_54_n78(net719_c1,net719);
INTERCONNECT SplitCLK_2_642_AND2T_46_n70(net720_c1,net720);
INTERCONNECT SplitCLK_4_641_AND2T_53_n77(net721_c1,net721);
INTERCONNECT SplitCLK_2_640_AND2T_61_n85(net722_c1,net722);
INTERCONNECT SplitCLK_4_639_AND2T_29_n53(net723_c1,net723);
INTERCONNECT SplitCLK_2_638_AND2T_28_n52(net724_c1,net724);
INTERCONNECT SplitCLK_2_637_AND2T_35_n59(net725_c1,net725);
INTERCONNECT SplitCLK_2_636_AND2T_51_n75(net726_c1,net726);
INTERCONNECT SplitCLK_2_635_AND2T_18_n42(net727_c1,net727);
INTERCONNECT SplitCLK_2_634_AND2T_25_n49(net728_c1,net728);
INTERCONNECT SplitCLK_4_633_AND2T_33_n57(net729_c1,net729);
INTERCONNECT SplitCLK_4_632_AND2T_32_n56(net730_c1,net730);
INTERCONNECT SplitCLK_4_631_AND2T_15_n39(net731_c1,net731);
INTERCONNECT SplitCLK_2_630_AND2T_22_n46(net732_c1,net732);
INTERCONNECT SplitCLK_4_629_AND2T_13_n37(net733_c1,net733);
INTERCONNECT SplitCLK_2_628_AND2T_21_n45(net734_c1,net734);
INTERCONNECT SplitCLK_2_627_AND2T_10_n34(net735_c1,net735);
INTERCONNECT SplitCLK_4_626_NOTT_8_n32(net736_c1,net736);
INTERCONNECT SplitCLK_2_625_AND2T_9_n33(net737_c1,net737);
INTERCONNECT SplitCLK_2_624_AND2T_139_n163(net738_c1,net738);
INTERCONNECT SplitCLK_2_623_AND2T_146_n182(net739_c1,net739);
INTERCONNECT SplitCLK_4_622_AND2T_129_n153(net740_c1,net740);
INTERCONNECT SplitCLK_2_621_AND2T_144_n180(net741_c1,net741);
INTERCONNECT SplitCLK_2_620_AND2T_128_n152(net742_c1,net742);
INTERCONNECT SplitCLK_2_619_AND2T_141_n177(net743_c1,net743);
INTERCONNECT SplitCLK_2_618_AND2T_133_n157(net744_c1,net744);
INTERCONNECT SplitCLK_4_617_AND2T_109_n133(net745_c1,net745);
INTERCONNECT SplitCLK_4_616_AND2T_140_n176(net746_c1,net746);
INTERCONNECT SplitCLK_4_615_AND2T_132_n156(net747_c1,net747);
INTERCONNECT SplitCLK_4_614_AND2T_123_n147(net748_c1,net748);
INTERCONNECT SplitCLK_4_613_AND2T_114_n138(net749_c1,net749);
INTERCONNECT SplitCLK_4_612_AND2T_122_n146(net750_c1,net750);
INTERCONNECT SplitCLK_2_611_AND2T_105_n129(net751_c1,net751);
INTERCONNECT SplitCLK_2_610_AND2T_113_n137(net752_c1,net752);
INTERCONNECT SplitCLK_4_609_AND2T_104_n128(net753_c1,net753);
INTERCONNECT SplitCLK_2_608_AND2T_103_n127(net754_c1,net754);
INTERCONNECT SplitCLK_2_607_AND2T_110_n134(net755_c1,net755);
INTERCONNECT SplitCLK_4_606_AND2T_101_n125(net756_c1,net756);
INTERCONNECT SplitCLK_4_605_XOR2T_55_n79(net757_c1,net757);
INTERCONNECT SplitCLK_4_604_XOR2T_45_n69(net758_c1,net758);
INTERCONNECT SplitCLK_2_603_XOR2T_36_n60(net759_c1,net759);
INTERCONNECT SplitCLK_4_602_DFFT_298__FPB_n754(net760_c1,net760);
INTERCONNECT SplitCLK_2_601_DFFT_288__FPB_n744(net761_c1,net761);
INTERCONNECT SplitCLK_2_600_DFFT_296__FPB_n752(net762_c1,net762);
INTERCONNECT SplitCLK_2_599_DFFT_199__FPB_n655(net763_c1,net763);
INTERCONNECT SplitCLK_4_598_DFFT_279__FPB_n735(net764_c1,net764);
INTERCONNECT SplitCLK_4_597_DFFT_287__FPB_n743(net765_c1,net765);
INTERCONNECT SplitCLK_2_596_SplitCLK_6_522(net766_c1,net766);
INTERCONNECT SplitCLK_2_596_SplitCLK_4_595(net767_c1,net767);
INTERCONNECT SplitCLK_4_595_SplitCLK_6_558(net768_c1,net768);
INTERCONNECT SplitCLK_4_595_SplitCLK_2_594(net769_c1,net769);
INTERCONNECT SplitCLK_2_594_SplitCLK_6_576(net770_c1,net770);
INTERCONNECT SplitCLK_2_594_SplitCLK_4_593(net771_c1,net771);
INTERCONNECT SplitCLK_4_593_SplitCLK_0_584(net772_c1,net772);
INTERCONNECT SplitCLK_4_593_SplitCLK_2_592(net773_c1,net773);
INTERCONNECT SplitCLK_2_592_SplitCLK_6_588(net774_c1,net774);
INTERCONNECT SplitCLK_2_592_SplitCLK_4_591(net775_c1,net775);
INTERCONNECT SplitCLK_4_591_SplitCLK_4_589(net776_c1,net776);
INTERCONNECT SplitCLK_4_591_SplitCLK_6_590(net777_c1,net777);
INTERCONNECT SplitCLK_6_590_SplitCLK_2_645(net778_c1,net778);
INTERCONNECT SplitCLK_6_590_SplitCLK_4_722(net779_c1,net779);
INTERCONNECT SplitCLK_4_589_SplitCLK_4_707(net780_c1,net780);
INTERCONNECT SplitCLK_4_589_SplitCLK_2_711(net781_c1,net781);
INTERCONNECT SplitCLK_6_588_SplitCLK_4_586(net782_c1,net782);
INTERCONNECT SplitCLK_6_588_SplitCLK_6_587(net783_c1,net783);
INTERCONNECT SplitCLK_6_587_SplitCLK_4_713(net784_c1,net784);
INTERCONNECT SplitCLK_6_587_SplitCLK_2_798(net785_c1,net785);
INTERCONNECT SplitCLK_4_586_SplitCLK_4_705(net786_c1,net786);
INTERCONNECT SplitCLK_4_586_SplitCLK_4_585(net787_c1,net787);
INTERCONNECT SplitCLK_4_585_AND2T_52_n76(net788_c1,net788);
INTERCONNECT SplitCLK_4_585_OR2T_77_n101(net789_c1,net789);
INTERCONNECT SplitCLK_0_584_SplitCLK_6_580(net790_c1,net790);
INTERCONNECT SplitCLK_0_584_SplitCLK_4_583(net791_c1,net791);
INTERCONNECT SplitCLK_4_583_SplitCLK_0_581(net792_c1,net792);
INTERCONNECT SplitCLK_4_583_SplitCLK_2_582(net793_c1,net793);
INTERCONNECT SplitCLK_2_582_SplitCLK_4_701(net794_c1,net794);
INTERCONNECT SplitCLK_2_582_SplitCLK_2_706(net795_c1,net795);
INTERCONNECT SplitCLK_0_581_SplitCLK_2_599(net796_c1,net796);
INTERCONNECT SplitCLK_0_581_SplitCLK_4_661(net797_c1,net797);
INTERCONNECT SplitCLK_6_580_SplitCLK_4_578(net798_c1,net798);
INTERCONNECT SplitCLK_6_580_SplitCLK_6_579(net799_c1,net799);
INTERCONNECT SplitCLK_6_579_SplitCLK_2_655(net800_c1,net800);
INTERCONNECT SplitCLK_6_579_SplitCLK_2_664(net801_c1,net801);
INTERCONNECT SplitCLK_4_578_SplitCLK_2_662(net802_c1,net802);
INTERCONNECT SplitCLK_4_578_SplitCLK_4_577(net803_c1,net803);
INTERCONNECT SplitCLK_4_577_AND2T_73_n97(net804_c1,net804);
INTERCONNECT SplitCLK_4_577_OR2T_37_n61(net805_c1,net805);
INTERCONNECT SplitCLK_6_576_SplitCLK_0_567(net806_c1,net806);
INTERCONNECT SplitCLK_6_576_SplitCLK_2_575(net807_c1,net807);
INTERCONNECT SplitCLK_2_575_SplitCLK_6_571(net808_c1,net808);
INTERCONNECT SplitCLK_2_575_SplitCLK_4_574(net809_c1,net809);
INTERCONNECT SplitCLK_4_574_SplitCLK_0_572(net810_c1,net810);
INTERCONNECT SplitCLK_4_574_SplitCLK_0_573(net811_c1,net811);
INTERCONNECT SplitCLK_0_573_SplitCLK_2_689(net812_c1,net812);
INTERCONNECT SplitCLK_0_573_SplitCLK_4_786(net813_c1,net813);
INTERCONNECT SplitCLK_0_572_SplitCLK_4_715(net814_c1,net814);
INTERCONNECT SplitCLK_0_572_SplitCLK_2_752(net815_c1,net815);
INTERCONNECT SplitCLK_6_571_SplitCLK_4_569(net816_c1,net816);
INTERCONNECT SplitCLK_6_571_SplitCLK_6_570(net817_c1,net817);
INTERCONNECT SplitCLK_6_570_SplitCLK_4_709(net818_c1,net818);
INTERCONNECT SplitCLK_6_570_SplitCLK_2_720(net819_c1,net819);
INTERCONNECT SplitCLK_4_569_SplitCLK_4_718(net820_c1,net820);
INTERCONNECT SplitCLK_4_569_SplitCLK_4_568(net821_c1,net821);
INTERCONNECT SplitCLK_4_568_AND2T_90_n114(net822_c1,net822);
INTERCONNECT SplitCLK_4_568_DFFT_223__FPB_n679(net823_c1,net823);
INTERCONNECT SplitCLK_0_567_SplitCLK_4_562(net824_c1,net824);
INTERCONNECT SplitCLK_0_567_SplitCLK_4_566(net825_c1,net825);
INTERCONNECT SplitCLK_4_566_SplitCLK_4_564(net826_c1,net826);
INTERCONNECT SplitCLK_4_566_SplitCLK_2_565(net827_c1,net827);
INTERCONNECT SplitCLK_2_565_SplitCLK_4_632(net828_c1,net828);
INTERCONNECT SplitCLK_2_565_SplitCLK_2_726(net829_c1,net829);
INTERCONNECT SplitCLK_4_564_SplitCLK_4_639(net830_c1,net830);
INTERCONNECT SplitCLK_4_564_SplitCLK_4_563(net831_c1,net831);
INTERCONNECT SplitCLK_4_563_DFFT_227__FPB_n683(net832_c1,net832);
INTERCONNECT SplitCLK_4_563_DFFT_228__FPB_n684(net833_c1,net833);
INTERCONNECT SplitCLK_4_562_SplitCLK_0_560(net834_c1,net834);
INTERCONNECT SplitCLK_4_562_SplitCLK_6_561(net835_c1,net835);
INTERCONNECT SplitCLK_6_561_SplitCLK_2_659(net836_c1,net836);
INTERCONNECT SplitCLK_6_561_SplitCLK_2_760(net837_c1,net837);
INTERCONNECT SplitCLK_0_560_SplitCLK_4_617(net838_c1,net838);
INTERCONNECT SplitCLK_0_560_SplitCLK_4_559(net839_c1,net839);
INTERCONNECT SplitCLK_4_559_AND2T_43_n67(net840_c1,net840);
INTERCONNECT SplitCLK_4_559_DFFT_205__FPB_n661(net841_c1,net841);
INTERCONNECT SplitCLK_6_558_SplitCLK_6_540(net842_c1,net842);
INTERCONNECT SplitCLK_6_558_SplitCLK_4_557(net843_c1,net843);
INTERCONNECT SplitCLK_4_557_SplitCLK_0_548(net844_c1,net844);
INTERCONNECT SplitCLK_4_557_SplitCLK_2_556(net845_c1,net845);
INTERCONNECT SplitCLK_2_556_SplitCLK_6_552(net846_c1,net846);
INTERCONNECT SplitCLK_2_556_SplitCLK_4_555(net847_c1,net847);
INTERCONNECT SplitCLK_4_555_SplitCLK_0_553(net848_c1,net848);
INTERCONNECT SplitCLK_4_555_SplitCLK_6_554(net849_c1,net849);
INTERCONNECT SplitCLK_6_554_SplitCLK_4_643(net850_c1,net850);
INTERCONNECT SplitCLK_6_554_SplitCLK_2_809(net851_c1,net851);
INTERCONNECT SplitCLK_0_553_SplitCLK_4_704(net852_c1,net852);
INTERCONNECT SplitCLK_0_553_SplitCLK_4_792(net853_c1,net853);
INTERCONNECT SplitCLK_6_552_SplitCLK_0_550(net854_c1,net854);
INTERCONNECT SplitCLK_6_552_SplitCLK_2_551(net855_c1,net855);
INTERCONNECT SplitCLK_2_551_SplitCLK_2_657(net856_c1,net856);
INTERCONNECT SplitCLK_2_551_SplitCLK_4_804(net857_c1,net857);
INTERCONNECT SplitCLK_0_550_SplitCLK_4_641(net858_c1,net858);
INTERCONNECT SplitCLK_0_550_SplitCLK_4_549(net859_c1,net859);
INTERCONNECT SplitCLK_4_549_DFFT_241__FPB_n697(net860_c1,net860);
INTERCONNECT SplitCLK_4_549_DFFT_189__FPB_n645(net861_c1,net861);
INTERCONNECT SplitCLK_0_548_SplitCLK_4_544(net862_c1,net862);
INTERCONNECT SplitCLK_0_548_SplitCLK_4_547(net863_c1,net863);
INTERCONNECT SplitCLK_4_547_SplitCLK_0_545(net864_c1,net864);
INTERCONNECT SplitCLK_4_547_SplitCLK_4_546(net865_c1,net865);
INTERCONNECT SplitCLK_4_546_SplitCLK_2_636(net866_c1,net866);
INTERCONNECT SplitCLK_4_546_SplitCLK_2_700(net867_c1,net867);
INTERCONNECT SplitCLK_0_545_SplitCLK_4_696(net868_c1,net868);
INTERCONNECT SplitCLK_0_545_SplitCLK_4_770(net869_c1,net869);
INTERCONNECT SplitCLK_4_544_SplitCLK_4_542(net870_c1,net870);
INTERCONNECT SplitCLK_4_544_SplitCLK_2_543(net871_c1,net871);
INTERCONNECT SplitCLK_2_543_SplitCLK_2_630(net872_c1,net872);
INTERCONNECT SplitCLK_2_543_SplitCLK_2_637(net873_c1,net873);
INTERCONNECT SplitCLK_4_542_SplitCLK_4_605(net874_c1,net874);
INTERCONNECT SplitCLK_4_542_SplitCLK_4_541(net875_c1,net875);
INTERCONNECT SplitCLK_4_541_OR2T_30_n54(net876_c1,net876);
INTERCONNECT SplitCLK_4_541_OR2T_23_n47(net877_c1,net877);
INTERCONNECT SplitCLK_6_540_SplitCLK_0_531(net878_c1,net878);
INTERCONNECT SplitCLK_6_540_SplitCLK_2_539(net879_c1,net879);
INTERCONNECT SplitCLK_2_539_SplitCLK_2_535(net880_c1,net880);
INTERCONNECT SplitCLK_2_539_SplitCLK_4_538(net881_c1,net881);
INTERCONNECT SplitCLK_4_538_SplitCLK_4_536(net882_c1,net882);
INTERCONNECT SplitCLK_4_538_SplitCLK_2_537(net883_c1,net883);
INTERCONNECT SplitCLK_2_537_SplitCLK_4_692(net884_c1,net884);
INTERCONNECT SplitCLK_2_537_SplitCLK_2_793(net885_c1,net885);
INTERCONNECT SplitCLK_4_536_SplitCLK_4_690(net886_c1,net886);
INTERCONNECT SplitCLK_4_536_SplitCLK_2_694(net887_c1,net887);
INTERCONNECT SplitCLK_2_535_SplitCLK_4_533(net888_c1,net888);
INTERCONNECT SplitCLK_2_535_SplitCLK_0_534(net889_c1,net889);
INTERCONNECT SplitCLK_0_534_SplitCLK_2_640(net890_c1,net890);
INTERCONNECT SplitCLK_0_534_SplitCLK_4_756(net891_c1,net891);
INTERCONNECT SplitCLK_4_533_SplitCLK_4_773(net892_c1,net892);
INTERCONNECT SplitCLK_4_533_SplitCLK_4_532(net893_c1,net893);
INTERCONNECT SplitCLK_4_532_OR2T_88_n112(net894_c1,net894);
INTERCONNECT SplitCLK_4_532_DFFT_190__FPB_n646(net895_c1,net895);
INTERCONNECT SplitCLK_0_531_SplitCLK_6_526(net896_c1,net896);
INTERCONNECT SplitCLK_0_531_SplitCLK_4_530(net897_c1,net897);
INTERCONNECT SplitCLK_4_530_SplitCLK_0_528(net898_c1,net898);
INTERCONNECT SplitCLK_4_530_SplitCLK_6_529(net899_c1,net899);
INTERCONNECT SplitCLK_6_529_SplitCLK_2_651(net900_c1,net900);
INTERCONNECT SplitCLK_6_529_SplitCLK_2_658(net901_c1,net901);
INTERCONNECT SplitCLK_0_528_SplitCLK_4_653(net902_c1,net902);
INTERCONNECT SplitCLK_0_528_SplitCLK_4_527(net903_c1,net903);
INTERCONNECT SplitCLK_4_527_AND2T_26_n50(net904_c1,net904);
INTERCONNECT SplitCLK_4_527_OR2T_69_n93(net905_c1,net905);
INTERCONNECT SplitCLK_6_526_SplitCLK_0_524(net906_c1,net906);
INTERCONNECT SplitCLK_6_526_SplitCLK_6_525(net907_c1,net907);
INTERCONNECT SplitCLK_6_525_SplitCLK_4_654(net908_c1,net908);
INTERCONNECT SplitCLK_6_525_SplitCLK_2_670(net909_c1,net909);
INTERCONNECT SplitCLK_0_524_SplitCLK_4_650(net910_c1,net910);
INTERCONNECT SplitCLK_0_524_SplitCLK_4_523(net911_c1,net911);
INTERCONNECT SplitCLK_4_523_AND2T_39_n63(net912_c1,net912);
INTERCONNECT SplitCLK_4_523_OR2T_111_n135(net913_c1,net913);
INTERCONNECT SplitCLK_6_522_SplitCLK_0_485(net914_c1,net914);
INTERCONNECT SplitCLK_6_522_SplitCLK_2_521(net915_c1,net915);
INTERCONNECT SplitCLK_2_521_SplitCLK_6_503(net916_c1,net916);
INTERCONNECT SplitCLK_2_521_SplitCLK_4_520(net917_c1,net917);
INTERCONNECT SplitCLK_4_520_SplitCLK_0_511(net918_c1,net918);
INTERCONNECT SplitCLK_4_520_SplitCLK_4_519(net919_c1,net919);
INTERCONNECT SplitCLK_4_519_SplitCLK_6_515(net920_c1,net920);
INTERCONNECT SplitCLK_4_519_SplitCLK_4_518(net921_c1,net921);
INTERCONNECT SplitCLK_4_518_SplitCLK_4_516(net922_c1,net922);
INTERCONNECT SplitCLK_4_518_SplitCLK_6_517(net923_c1,net923);
INTERCONNECT SplitCLK_6_517_SplitCLK_2_716(net924_c1,net924);
INTERCONNECT SplitCLK_6_517_SplitCLK_4_728(net925_c1,net925);
INTERCONNECT SplitCLK_4_516_SplitCLK_4_724(net926_c1,net926);
INTERCONNECT SplitCLK_4_516_SplitCLK_2_736(net927_c1,net927);
INTERCONNECT SplitCLK_6_515_SplitCLK_4_513(net928_c1,net928);
INTERCONNECT SplitCLK_6_515_SplitCLK_6_514(net929_c1,net929);
INTERCONNECT SplitCLK_6_514_SplitCLK_2_687(net930_c1,net930);
INTERCONNECT SplitCLK_6_514_SplitCLK_4_758(net931_c1,net931);
INTERCONNECT SplitCLK_4_513_SplitCLK_4_725(net932_c1,net932);
INTERCONNECT SplitCLK_4_513_SplitCLK_4_512(net933_c1,net933);
INTERCONNECT SplitCLK_4_512_NOTT_149_n197(net934_c1,net934);
INTERCONNECT SplitCLK_4_512_DFFT_184__FPB_n640(net935_c1,net935);
INTERCONNECT SplitCLK_0_511_SplitCLK_6_507(net936_c1,net936);
INTERCONNECT SplitCLK_0_511_SplitCLK_4_510(net937_c1,net937);
INTERCONNECT SplitCLK_4_510_SplitCLK_0_508(net938_c1,net938);
INTERCONNECT SplitCLK_4_510_SplitCLK_6_509(net939_c1,net939);
INTERCONNECT SplitCLK_6_509_SplitCLK_2_688(net940_c1,net940);
INTERCONNECT SplitCLK_6_509_SplitCLK_4_723(net941_c1,net941);
INTERCONNECT SplitCLK_0_508_SplitCLK_4_668(net942_c1,net942);
INTERCONNECT SplitCLK_0_508_SplitCLK_4_795(net943_c1,net943);
INTERCONNECT SplitCLK_6_507_SplitCLK_4_505(net944_c1,net944);
INTERCONNECT SplitCLK_6_507_SplitCLK_4_506(net945_c1,net945);
INTERCONNECT SplitCLK_4_506_SplitCLK_2_667(net946_c1,net946);
INTERCONNECT SplitCLK_4_506_SplitCLK_2_767(net947_c1,net947);
INTERCONNECT SplitCLK_4_505_SplitCLK_4_616(net948_c1,net948);
INTERCONNECT SplitCLK_4_505_SplitCLK_4_504(net949_c1,net949);
INTERCONNECT SplitCLK_4_504_DFFT_220__FPB_n676(net950_c1,net950);
INTERCONNECT SplitCLK_4_504_DFFT_167__FBL_n623(net951_c1,net951);
INTERCONNECT SplitCLK_6_503_SplitCLK_0_494(net952_c1,net952);
INTERCONNECT SplitCLK_6_503_SplitCLK_2_502(net953_c1,net953);
INTERCONNECT SplitCLK_2_502_SplitCLK_0_498(net954_c1,net954);
INTERCONNECT SplitCLK_2_502_SplitCLK_4_501(net955_c1,net955);
INTERCONNECT SplitCLK_4_501_SplitCLK_4_499(net956_c1,net956);
INTERCONNECT SplitCLK_4_501_SplitCLK_6_500(net957_c1,net957);
INTERCONNECT SplitCLK_6_500_SplitCLK_4_710(net958_c1,net958);
INTERCONNECT SplitCLK_6_500_SplitCLK_2_775(net959_c1,net959);
INTERCONNECT SplitCLK_4_499_SplitCLK_2_721(net960_c1,net960);
INTERCONNECT SplitCLK_4_499_SplitCLK_4_729(net961_c1,net961);
INTERCONNECT SplitCLK_0_498_SplitCLK_0_496(net962_c1,net962);
INTERCONNECT SplitCLK_0_498_SplitCLK_2_497(net963_c1,net963);
INTERCONNECT SplitCLK_2_497_SplitCLK_4_598(net964_c1,net964);
INTERCONNECT SplitCLK_2_497_SplitCLK_2_665(net965_c1,net965);
INTERCONNECT SplitCLK_0_496_SplitCLK_4_698(net966_c1,net966);
INTERCONNECT SplitCLK_0_496_SplitCLK_0_495(net967_c1,net967);
INTERCONNECT SplitCLK_0_495_DFFT_283__FPB_n739(net968_c1,net968);
INTERCONNECT SplitCLK_0_495_DFFT_284__FPB_n740(net969_c1,net969);
INTERCONNECT SplitCLK_0_494_SplitCLK_6_489(net970_c1,net970);
INTERCONNECT SplitCLK_0_494_SplitCLK_4_493(net971_c1,net971);
INTERCONNECT SplitCLK_4_493_SplitCLK_2_491(net972_c1,net972);
INTERCONNECT SplitCLK_4_493_SplitCLK_6_492(net973_c1,net973);
INTERCONNECT SplitCLK_6_492_SplitCLK_2_625(net974_c1,net974);
INTERCONNECT SplitCLK_6_492_SplitCLK_4_737(net975_c1,net975);
INTERCONNECT SplitCLK_2_491_SplitCLK_2_741(net976_c1,net976);
INTERCONNECT SplitCLK_2_491_SplitCLK_4_490(net977_c1,net977);
INTERCONNECT SplitCLK_4_490_DFFT_221__FPB_n677(net978_c1,net978);
INTERCONNECT SplitCLK_4_490_DFFT_174__FPB_n630(net979_c1,net979);
INTERCONNECT SplitCLK_6_489_SplitCLK_0_487(net980_c1,net980);
INTERCONNECT SplitCLK_6_489_SplitCLK_6_488(net981_c1,net981);
INTERCONNECT SplitCLK_6_488_SplitCLK_4_781(net982_c1,net982);
INTERCONNECT SplitCLK_6_488_SplitCLK_2_788(net983_c1,net983);
INTERCONNECT SplitCLK_0_487_SplitCLK_4_750(net984_c1,net984);
INTERCONNECT SplitCLK_0_487_SplitCLK_4_486(net985_c1,net985);
INTERCONNECT SplitCLK_4_486_DFFT_292_state_obs1(net986_c1,net986);
INTERCONNECT SplitCLK_4_486_DFFT_291__FPB_n747(net987_c1,net987);
INTERCONNECT SplitCLK_0_485_SplitCLK_6_466(net988_c1,net988);
INTERCONNECT SplitCLK_0_485_SplitCLK_4_484(net989_c1,net989);
INTERCONNECT SplitCLK_4_484_SplitCLK_0_475(net990_c1,net990);
INTERCONNECT SplitCLK_4_484_SplitCLK_2_483(net991_c1,net991);
INTERCONNECT SplitCLK_2_483_SplitCLK_6_479(net992_c1,net992);
INTERCONNECT SplitCLK_2_483_SplitCLK_2_482(net993_c1,net993);
INTERCONNECT SplitCLK_2_482_SplitCLK_0_480(net994_c1,net994);
INTERCONNECT SplitCLK_2_482_SplitCLK_6_481(net995_c1,net995);
INTERCONNECT SplitCLK_6_481_SplitCLK_2_635(net996_c1,net996);
INTERCONNECT SplitCLK_6_481_SplitCLK_2_642(net997_c1,net997);
INTERCONNECT SplitCLK_0_480_SplitCLK_4_674(net998_c1,net998);
INTERCONNECT SplitCLK_0_480_SplitCLK_4_785(net999_c1,net999);
INTERCONNECT SplitCLK_6_479_SplitCLK_4_477(net1000_c1,net1000);
INTERCONNECT SplitCLK_6_479_SplitCLK_6_478(net1001_c1,net1001);
INTERCONNECT SplitCLK_6_478_SplitCLK_2_739(net1002_c1,net1002);
INTERCONNECT SplitCLK_6_478_SplitCLK_4_742(net1003_c1,net1003);
INTERCONNECT SplitCLK_4_477_SplitCLK_4_763(net1004_c1,net1004);
INTERCONNECT SplitCLK_4_477_SplitCLK_4_476(net1005_c1,net1005);
INTERCONNECT SplitCLK_4_476_AND2T_98_n122(net1006_c1,net1006);
INTERCONNECT SplitCLK_4_476_DFFT_160__FBL_n616(net1007_c1,net1007);
INTERCONNECT SplitCLK_0_475_SplitCLK_6_470(net1008_c1,net1008);
INTERCONNECT SplitCLK_0_475_SplitCLK_4_474(net1009_c1,net1009);
INTERCONNECT SplitCLK_4_474_SplitCLK_4_472(net1010_c1,net1010);
INTERCONNECT SplitCLK_4_474_SplitCLK_2_473(net1011_c1,net1011);
INTERCONNECT SplitCLK_2_473_SplitCLK_2_646(net1012_c1,net1012);
INTERCONNECT SplitCLK_2_473_SplitCLK_2_777(net1013_c1,net1013);
INTERCONNECT SplitCLK_4_472_SplitCLK_4_673(net1014_c1,net1014);
INTERCONNECT SplitCLK_4_472_SplitCLK_4_471(net1015_c1,net1015);
INTERCONNECT SplitCLK_4_471_AND2T_44_n68(net1016_c1,net1016);
INTERCONNECT SplitCLK_4_471_DFFT_240__FPB_n696(net1017_c1,net1017);
INTERCONNECT SplitCLK_6_470_SplitCLK_0_468(net1018_c1,net1018);
INTERCONNECT SplitCLK_6_470_SplitCLK_6_469(net1019_c1,net1019);
INTERCONNECT SplitCLK_6_469_SplitCLK_2_634(net1020_c1,net1020);
INTERCONNECT SplitCLK_6_469_SplitCLK_2_808(net1021_c1,net1021);
INTERCONNECT SplitCLK_0_468_SplitCLK_4_730(net1022_c1,net1022);
INTERCONNECT SplitCLK_0_468_SplitCLK_4_467(net1023_c1,net1023);
INTERCONNECT SplitCLK_4_467_AND2T_143_n179(net1024_c1,net1024);
INTERCONNECT SplitCLK_4_467_AND2T_145_n181(net1025_c1,net1025);
INTERCONNECT SplitCLK_6_466_SplitCLK_4_457(net1026_c1,net1026);
INTERCONNECT SplitCLK_6_466_SplitCLK_6_465(net1027_c1,net1027);
INTERCONNECT SplitCLK_6_465_SplitCLK_6_461(net1028_c1,net1028);
INTERCONNECT SplitCLK_6_465_SplitCLK_4_464(net1029_c1,net1029);
INTERCONNECT SplitCLK_4_464_SplitCLK_4_462(net1030_c1,net1030);
INTERCONNECT SplitCLK_4_464_SplitCLK_2_463(net1031_c1,net1031);
INTERCONNECT SplitCLK_2_463_SplitCLK_2_702(net1032_c1,net1032);
INTERCONNECT SplitCLK_2_463_SplitCLK_4_765(net1033_c1,net1033);
INTERCONNECT SplitCLK_4_462_SplitCLK_4_751(net1034_c1,net1034);
INTERCONNECT SplitCLK_4_462_SplitCLK_2_757(net1035_c1,net1035);
INTERCONNECT SplitCLK_6_461_SplitCLK_0_459(net1036_c1,net1036);
INTERCONNECT SplitCLK_6_461_SplitCLK_2_460(net1037_c1,net1037);
INTERCONNECT SplitCLK_2_460_SplitCLK_2_601(net1038_c1,net1038);
INTERCONNECT SplitCLK_2_460_SplitCLK_4_807(net1039_c1,net1039);
INTERCONNECT SplitCLK_0_459_SplitCLK_4_597(net1040_c1,net1040);
INTERCONNECT SplitCLK_0_459_SplitCLK_4_458(net1041_c1,net1041);
INTERCONNECT SplitCLK_4_458_DFFT_289__FPB_n745(net1042_c1,net1042);
INTERCONNECT SplitCLK_4_458_DFFT_290__FPB_n746(net1043_c1,net1043);
INTERCONNECT SplitCLK_4_457_SplitCLK_0_452(net1044_c1,net1044);
INTERCONNECT SplitCLK_4_457_SplitCLK_4_456(net1045_c1,net1045);
INTERCONNECT SplitCLK_4_456_SplitCLK_0_454(net1046_c1,net1046);
INTERCONNECT SplitCLK_4_456_SplitCLK_6_455(net1047_c1,net1047);
INTERCONNECT SplitCLK_6_455_SplitCLK_2_627(net1048_c1,net1048);
INTERCONNECT SplitCLK_6_455_SplitCLK_4_747(net1049_c1,net1049);
INTERCONNECT SplitCLK_0_454_SplitCLK_4_666(net1050_c1,net1050);
INTERCONNECT SplitCLK_0_454_SplitCLK_4_453(net1051_c1,net1051);
INTERCONNECT SplitCLK_4_453_DFFT_234__FPB_n690(net1052_c1,net1052);
INTERCONNECT SplitCLK_4_453_DFFT_235__FPB_n691(net1053_c1,net1053);
INTERCONNECT SplitCLK_0_452_SplitCLK_4_450(net1054_c1,net1054);
INTERCONNECT SplitCLK_0_452_SplitCLK_6_451(net1055_c1,net1055);
INTERCONNECT SplitCLK_6_451_SplitCLK_4_602(net1056_c1,net1056);
INTERCONNECT SplitCLK_6_451_SplitCLK_2_686(net1057_c1,net1057);
INTERCONNECT SplitCLK_4_450_SplitCLK_2_774(net1058_c1,net1058);
INTERCONNECT SplitCLK_4_450_SplitCLK_4_449(net1059_c1,net1059);
INTERCONNECT SplitCLK_4_449_DFFT_297__FPB_n753(net1060_c1,net1060);
INTERCONNECT SplitCLK_4_449_DFFT_175__FPB_n631(net1061_c1,net1061);
INTERCONNECT SplitCLK_0_448_SplitCLK_6_373(net1062_c1,net1062);
INTERCONNECT SplitCLK_0_448_SplitCLK_4_447(net1063_c1,net1063);
INTERCONNECT SplitCLK_4_447_SplitCLK_0_410(net1064_c1,net1064);
INTERCONNECT SplitCLK_4_447_SplitCLK_2_446(net1065_c1,net1065);
INTERCONNECT SplitCLK_2_446_SplitCLK_6_428(net1066_c1,net1066);
INTERCONNECT SplitCLK_2_446_SplitCLK_4_445(net1067_c1,net1067);
INTERCONNECT SplitCLK_4_445_SplitCLK_0_436(net1068_c1,net1068);
INTERCONNECT SplitCLK_4_445_SplitCLK_6_444(net1069_c1,net1069);
INTERCONNECT SplitCLK_6_444_SplitCLK_0_440(net1070_c1,net1070);
INTERCONNECT SplitCLK_6_444_SplitCLK_2_443(net1071_c1,net1071);
INTERCONNECT SplitCLK_2_443_SplitCLK_4_441(net1072_c1,net1072);
INTERCONNECT SplitCLK_2_443_SplitCLK_2_442(net1073_c1,net1073);
INTERCONNECT SplitCLK_2_442_SplitCLK_2_649(net1074_c1,net1074);
INTERCONNECT SplitCLK_2_442_SplitCLK_4_771(net1075_c1,net1075);
INTERCONNECT SplitCLK_4_441_SplitCLK_4_784(net1076_c1,net1076);
INTERCONNECT SplitCLK_4_441_SplitCLK_2_789(net1077_c1,net1077);
INTERCONNECT SplitCLK_0_440_SplitCLK_4_438(net1078_c1,net1078);
INTERCONNECT SplitCLK_0_440_SplitCLK_6_439(net1079_c1,net1079);
INTERCONNECT SplitCLK_6_439_SplitCLK_4_647(net1080_c1,net1080);
INTERCONNECT SplitCLK_6_439_SplitCLK_2_717(net1081_c1,net1081);
INTERCONNECT SplitCLK_4_438_SplitCLK_2_697(net1082_c1,net1082);
INTERCONNECT SplitCLK_4_438_SplitCLK_4_437(net1083_c1,net1083);
INTERCONNECT SplitCLK_4_437_AND2T_56_n80(net1084_c1,net1084);
INTERCONNECT SplitCLK_4_437_DFFT_211__FPB_n667(net1085_c1,net1085);
INTERCONNECT SplitCLK_0_436_SplitCLK_6_432(net1086_c1,net1086);
INTERCONNECT SplitCLK_0_436_SplitCLK_4_435(net1087_c1,net1087);
INTERCONNECT SplitCLK_4_435_SplitCLK_4_433(net1088_c1,net1088);
INTERCONNECT SplitCLK_4_435_SplitCLK_6_434(net1089_c1,net1089);
INTERCONNECT SplitCLK_6_434_SplitCLK_4_776(net1090_c1,net1090);
INTERCONNECT SplitCLK_6_434_SplitCLK_2_782(net1091_c1,net1091);
INTERCONNECT SplitCLK_4_433_SplitCLK_4_734(net1092_c1,net1092);
INTERCONNECT SplitCLK_4_433_SplitCLK_2_761(net1093_c1,net1093);
INTERCONNECT SplitCLK_6_432_SplitCLK_0_430(net1094_c1,net1094);
INTERCONNECT SplitCLK_6_432_SplitCLK_4_431(net1095_c1,net1095);
INTERCONNECT SplitCLK_4_431_SplitCLK_2_663(net1096_c1,net1096);
INTERCONNECT SplitCLK_4_431_SplitCLK_2_712(net1097_c1,net1097);
INTERCONNECT SplitCLK_0_430_SplitCLK_4_656(net1098_c1,net1098);
INTERCONNECT SplitCLK_0_430_SplitCLK_4_429(net1099_c1,net1099);
INTERCONNECT SplitCLK_4_429_AND2T_106_n130(net1100_c1,net1100);
INTERCONNECT SplitCLK_4_429_DFFT_245__FPB_n701(net1101_c1,net1101);
INTERCONNECT SplitCLK_6_428_SplitCLK_0_419(net1102_c1,net1102);
INTERCONNECT SplitCLK_6_428_SplitCLK_2_427(net1103_c1,net1103);
INTERCONNECT SplitCLK_2_427_SplitCLK_6_423(net1104_c1,net1104);
INTERCONNECT SplitCLK_2_427_SplitCLK_0_426(net1105_c1,net1105);
INTERCONNECT SplitCLK_0_426_SplitCLK_0_424(net1106_c1,net1106);
INTERCONNECT SplitCLK_0_426_SplitCLK_2_425(net1107_c1,net1107);
INTERCONNECT SplitCLK_2_425_SplitCLK_2_660(net1108_c1,net1108);
INTERCONNECT SplitCLK_2_425_SplitCLK_4_675(net1109_c1,net1109);
INTERCONNECT SplitCLK_0_424_SplitCLK_4_606(net1110_c1,net1110);
INTERCONNECT SplitCLK_0_424_SplitCLK_4_633(net1111_c1,net1111);
INTERCONNECT SplitCLK_6_423_SplitCLK_0_421(net1112_c1,net1112);
INTERCONNECT SplitCLK_6_423_SplitCLK_6_422(net1113_c1,net1113);
INTERCONNECT SplitCLK_6_422_SplitCLK_2_644(net1114_c1,net1114);
INTERCONNECT SplitCLK_6_422_SplitCLK_4_676(net1115_c1,net1115);
INTERCONNECT SplitCLK_0_421_SplitCLK_4_652(net1116_c1,net1116);
INTERCONNECT SplitCLK_0_421_SplitCLK_4_420(net1117_c1,net1117);
INTERCONNECT SplitCLK_4_420_OR2T_130_n154(net1118_c1,net1118);
INTERCONNECT SplitCLK_4_420_AND2T_86_n110(net1119_c1,net1119);
INTERCONNECT SplitCLK_0_419_SplitCLK_4_414(net1120_c1,net1120);
INTERCONNECT SplitCLK_0_419_SplitCLK_4_418(net1121_c1,net1121);
INTERCONNECT SplitCLK_4_418_SplitCLK_4_416(net1122_c1,net1122);
INTERCONNECT SplitCLK_4_418_SplitCLK_2_417(net1123_c1,net1123);
INTERCONNECT SplitCLK_2_417_SplitCLK_2_671(net1124_c1,net1124);
INTERCONNECT SplitCLK_2_417_SplitCLK_4_691(net1125_c1,net1125);
INTERCONNECT SplitCLK_4_416_SplitCLK_4_615(net1126_c1,net1126);
INTERCONNECT SplitCLK_4_416_SplitCLK_4_415(net1127_c1,net1127);
INTERCONNECT SplitCLK_4_415_OR2T_134_n158(net1128_c1,net1128);
INTERCONNECT SplitCLK_4_415_DFFT_264__FPB_n720(net1129_c1,net1129);
INTERCONNECT SplitCLK_4_414_SplitCLK_4_412(net1130_c1,net1130);
INTERCONNECT SplitCLK_4_414_SplitCLK_2_413(net1131_c1,net1131);
INTERCONNECT SplitCLK_2_413_SplitCLK_2_607(net1132_c1,net1132);
INTERCONNECT SplitCLK_2_413_SplitCLK_2_681(net1133_c1,net1133);
INTERCONNECT SplitCLK_4_412_SplitCLK_2_608(net1134_c1,net1134);
INTERCONNECT SplitCLK_4_412_SplitCLK_4_411(net1135_c1,net1135);
INTERCONNECT SplitCLK_4_411_AND2T_16_n40(net1136_c1,net1136);
INTERCONNECT SplitCLK_4_411_OR2T_131_n155(net1137_c1,net1137);
INTERCONNECT SplitCLK_0_410_SplitCLK_6_391(net1138_c1,net1138);
INTERCONNECT SplitCLK_0_410_SplitCLK_4_409(net1139_c1,net1139);
INTERCONNECT SplitCLK_4_409_SplitCLK_0_400(net1140_c1,net1140);
INTERCONNECT SplitCLK_4_409_SplitCLK_2_408(net1141_c1,net1141);
INTERCONNECT SplitCLK_2_408_SplitCLK_6_404(net1142_c1,net1142);
INTERCONNECT SplitCLK_2_408_SplitCLK_4_407(net1143_c1,net1143);
INTERCONNECT SplitCLK_4_407_SplitCLK_4_405(net1144_c1,net1144);
INTERCONNECT SplitCLK_4_407_SplitCLK_6_406(net1145_c1,net1145);
INTERCONNECT SplitCLK_6_406_SplitCLK_4_699(net1146_c1,net1146);
INTERCONNECT SplitCLK_6_406_SplitCLK_2_703(net1147_c1,net1147);
INTERCONNECT SplitCLK_4_405_SplitCLK_2_769(net1148_c1,net1148);
INTERCONNECT SplitCLK_4_405_SplitCLK_4_797(net1149_c1,net1149);
INTERCONNECT SplitCLK_6_404_SplitCLK_4_402(net1150_c1,net1150);
INTERCONNECT SplitCLK_6_404_SplitCLK_6_403(net1151_c1,net1151);
INTERCONNECT SplitCLK_6_403_SplitCLK_4_609(net1152_c1,net1152);
INTERCONNECT SplitCLK_6_403_SplitCLK_2_618(net1153_c1,net1153);
INTERCONNECT SplitCLK_4_402_SplitCLK_4_708(net1154_c1,net1154);
INTERCONNECT SplitCLK_4_402_SplitCLK_4_401(net1155_c1,net1155);
INTERCONNECT SplitCLK_4_401_OR2T_107_n131(net1156_c1,net1156);
INTERCONNECT SplitCLK_4_401_DFFT_153__FPB_n207(net1157_c1,net1157);
INTERCONNECT SplitCLK_0_400_SplitCLK_0_395(net1158_c1,net1158);
INTERCONNECT SplitCLK_0_400_SplitCLK_4_399(net1159_c1,net1159);
INTERCONNECT SplitCLK_4_399_SplitCLK_4_397(net1160_c1,net1160);
INTERCONNECT SplitCLK_4_399_SplitCLK_4_398(net1161_c1,net1161);
INTERCONNECT SplitCLK_4_398_SplitCLK_4_755(net1162_c1,net1162);
INTERCONNECT SplitCLK_4_398_SplitCLK_2_803(net1163_c1,net1163);
INTERCONNECT SplitCLK_4_397_SplitCLK_2_738(net1164_c1,net1164);
INTERCONNECT SplitCLK_4_397_SplitCLK_4_396(net1165_c1,net1165);
INTERCONNECT SplitCLK_4_396_DFFT_243__FPB_n699(net1166_c1,net1166);
INTERCONNECT SplitCLK_4_396_DFFT_265__FPB_n721(net1167_c1,net1167);
INTERCONNECT SplitCLK_0_395_SplitCLK_0_393(net1168_c1,net1168);
INTERCONNECT SplitCLK_0_395_SplitCLK_6_394(net1169_c1,net1169);
INTERCONNECT SplitCLK_6_394_SplitCLK_2_611(net1170_c1,net1170);
INTERCONNECT SplitCLK_6_394_SplitCLK_4_743(net1171_c1,net1171);
INTERCONNECT SplitCLK_0_393_SplitCLK_4_778(net1172_c1,net1172);
INTERCONNECT SplitCLK_0_393_SplitCLK_0_392(net1173_c1,net1173);
INTERCONNECT SplitCLK_0_392_DFFT_266__FPB_n722(net1174_c1,net1174);
INTERCONNECT SplitCLK_0_392_DFFT_258__FPB_n714(net1175_c1,net1175);
INTERCONNECT SplitCLK_6_391_SplitCLK_4_382(net1176_c1,net1176);
INTERCONNECT SplitCLK_6_391_SplitCLK_2_390(net1177_c1,net1177);
INTERCONNECT SplitCLK_2_390_SplitCLK_6_386(net1178_c1,net1178);
INTERCONNECT SplitCLK_2_390_SplitCLK_4_389(net1179_c1,net1179);
INTERCONNECT SplitCLK_4_389_SplitCLK_0_387(net1180_c1,net1180);
INTERCONNECT SplitCLK_4_389_SplitCLK_4_388(net1181_c1,net1181);
INTERCONNECT SplitCLK_4_388_SplitCLK_2_603(net1182_c1,net1182);
INTERCONNECT SplitCLK_4_388_SplitCLK_4_799(net1183_c1,net1183);
INTERCONNECT SplitCLK_0_387_SplitCLK_2_754(net1184_c1,net1184);
INTERCONNECT SplitCLK_0_387_SplitCLK_4_791(net1185_c1,net1185);
INTERCONNECT SplitCLK_6_386_SplitCLK_2_384(net1186_c1,net1186);
INTERCONNECT SplitCLK_6_386_SplitCLK_6_385(net1187_c1,net1187);
INTERCONNECT SplitCLK_6_385_SplitCLK_2_610(net1188_c1,net1188);
INTERCONNECT SplitCLK_6_385_SplitCLK_2_683(net1189_c1,net1189);
INTERCONNECT SplitCLK_2_384_SplitCLK_2_678(net1190_c1,net1190);
INTERCONNECT SplitCLK_2_384_SplitCLK_4_383(net1191_c1,net1191);
INTERCONNECT SplitCLK_4_383_OR2T_115_n139(net1192_c1,net1192);
INTERCONNECT SplitCLK_4_383_OR2T_116_n140(net1193_c1,net1193);
INTERCONNECT SplitCLK_4_382_SplitCLK_6_377(net1194_c1,net1194);
INTERCONNECT SplitCLK_4_382_SplitCLK_6_381(net1195_c1,net1195);
INTERCONNECT SplitCLK_6_381_SplitCLK_0_379(net1196_c1,net1196);
INTERCONNECT SplitCLK_6_381_SplitCLK_2_380(net1197_c1,net1197);
INTERCONNECT SplitCLK_2_380_SplitCLK_2_677(net1198_c1,net1198);
INTERCONNECT SplitCLK_2_380_SplitCLK_4_744(net1199_c1,net1199);
INTERCONNECT SplitCLK_0_379_SplitCLK_4_614(net1200_c1,net1200);
INTERCONNECT SplitCLK_0_379_SplitCLK_4_378(net1201_c1,net1201);
INTERCONNECT SplitCLK_4_378_DFFT_261__FPB_n717(net1202_c1,net1202);
INTERCONNECT SplitCLK_4_378_DFFT_262__FPB_n718(net1203_c1,net1203);
INTERCONNECT SplitCLK_6_377_SplitCLK_4_375(net1204_c1,net1204);
INTERCONNECT SplitCLK_6_377_SplitCLK_6_376(net1205_c1,net1205);
INTERCONNECT SplitCLK_6_376_SplitCLK_2_680(net1206_c1,net1206);
INTERCONNECT SplitCLK_6_376_SplitCLK_4_684(net1207_c1,net1207);
INTERCONNECT SplitCLK_4_375_SplitCLK_4_612(net1208_c1,net1208);
INTERCONNECT SplitCLK_4_375_SplitCLK_4_374(net1209_c1,net1209);
INTERCONNECT SplitCLK_4_374_AND2T_124_n148(net1210_c1,net1210);
INTERCONNECT SplitCLK_4_374_OR2T_126_n150(net1211_c1,net1211);
INTERCONNECT SplitCLK_6_373_SplitCLK_0_336(net1212_c1,net1212);
INTERCONNECT SplitCLK_6_373_SplitCLK_6_372(net1213_c1,net1213);
INTERCONNECT SplitCLK_6_372_SplitCLK_6_354(net1214_c1,net1214);
INTERCONNECT SplitCLK_6_372_SplitCLK_4_371(net1215_c1,net1215);
INTERCONNECT SplitCLK_4_371_SplitCLK_0_362(net1216_c1,net1216);
INTERCONNECT SplitCLK_4_371_SplitCLK_4_370(net1217_c1,net1217);
INTERCONNECT SplitCLK_4_370_SplitCLK_6_366(net1218_c1,net1218);
INTERCONNECT SplitCLK_4_370_SplitCLK_4_369(net1219_c1,net1219);
INTERCONNECT SplitCLK_4_369_SplitCLK_4_367(net1220_c1,net1220);
INTERCONNECT SplitCLK_4_369_SplitCLK_2_368(net1221_c1,net1221);
INTERCONNECT SplitCLK_2_368_SplitCLK_2_620(net1222_c1,net1222);
INTERCONNECT SplitCLK_2_368_SplitCLK_2_648(net1223_c1,net1223);
INTERCONNECT SplitCLK_4_367_SplitCLK_2_621(net1224_c1,net1224);
INTERCONNECT SplitCLK_4_367_SplitCLK_4_802(net1225_c1,net1225);
INTERCONNECT SplitCLK_6_366_SplitCLK_4_364(net1226_c1,net1226);
INTERCONNECT SplitCLK_6_366_SplitCLK_2_365(net1227_c1,net1227);
INTERCONNECT SplitCLK_2_365_SplitCLK_2_695(net1228_c1,net1228);
INTERCONNECT SplitCLK_2_365_SplitCLK_2_762(net1229_c1,net1229);
INTERCONNECT SplitCLK_4_364_SplitCLK_4_604(net1230_c1,net1230);
INTERCONNECT SplitCLK_4_364_SplitCLK_4_363(net1231_c1,net1231);
INTERCONNECT SplitCLK_4_363_AND2T_24_n48(net1232_c1,net1232);
INTERCONNECT SplitCLK_4_363_OR2T_100_n124(net1233_c1,net1233);
INTERCONNECT SplitCLK_0_362_SplitCLK_4_358(net1234_c1,net1234);
INTERCONNECT SplitCLK_0_362_SplitCLK_4_361(net1235_c1,net1235);
INTERCONNECT SplitCLK_4_361_SplitCLK_0_359(net1236_c1,net1236);
INTERCONNECT SplitCLK_4_361_SplitCLK_4_360(net1237_c1,net1237);
INTERCONNECT SplitCLK_4_360_SplitCLK_2_623(net1238_c1,net1238);
INTERCONNECT SplitCLK_4_360_SplitCLK_2_693(net1239_c1,net1239);
INTERCONNECT SplitCLK_0_359_SplitCLK_4_622(net1240_c1,net1240);
INTERCONNECT SplitCLK_0_359_SplitCLK_4_753(net1241_c1,net1241);
INTERCONNECT SplitCLK_4_358_SplitCLK_0_356(net1242_c1,net1242);
INTERCONNECT SplitCLK_4_358_SplitCLK_2_357(net1243_c1,net1243);
INTERCONNECT SplitCLK_2_357_SplitCLK_2_638(net1244_c1,net1244);
INTERCONNECT SplitCLK_2_357_SplitCLK_4_783(net1245_c1,net1245);
INTERCONNECT SplitCLK_0_356_SplitCLK_4_669(net1246_c1,net1246);
INTERCONNECT SplitCLK_0_356_SplitCLK_4_355(net1247_c1,net1247);
INTERCONNECT SplitCLK_4_355_AND2T_27_n51(net1248_c1,net1248);
INTERCONNECT SplitCLK_4_355_DFFT_171__FBL_n627(net1249_c1,net1249);
INTERCONNECT SplitCLK_6_354_SplitCLK_6_345(net1250_c1,net1250);
INTERCONNECT SplitCLK_6_354_SplitCLK_6_353(net1251_c1,net1251);
INTERCONNECT SplitCLK_6_353_SplitCLK_6_349(net1252_c1,net1252);
INTERCONNECT SplitCLK_6_353_SplitCLK_4_352(net1253_c1,net1253);
INTERCONNECT SplitCLK_4_352_SplitCLK_0_350(net1254_c1,net1254);
INTERCONNECT SplitCLK_4_352_SplitCLK_2_351(net1255_c1,net1255);
INTERCONNECT SplitCLK_2_351_SplitCLK_4_629(net1256_c1,net1256);
INTERCONNECT SplitCLK_2_351_SplitCLK_2_731(net1257_c1,net1257);
INTERCONNECT SplitCLK_0_350_SplitCLK_4_672(net1258_c1,net1258);
INTERCONNECT SplitCLK_0_350_SplitCLK_2_800(net1259_c1,net1259);
INTERCONNECT SplitCLK_6_349_SplitCLK_0_347(net1260_c1,net1260);
INTERCONNECT SplitCLK_6_349_SplitCLK_2_348(net1261_c1,net1261);
INTERCONNECT SplitCLK_2_348_SplitCLK_2_600(net1262_c1,net1262);
INTERCONNECT SplitCLK_2_348_SplitCLK_4_626(net1263_c1,net1263);
INTERCONNECT SplitCLK_0_347_SplitCLK_4_746(net1264_c1,net1264);
INTERCONNECT SplitCLK_0_347_SplitCLK_0_346(net1265_c1,net1265);
INTERCONNECT SplitCLK_0_346_DFFT_295__FPB_n751(net1266_c1,net1266);
INTERCONNECT SplitCLK_0_346_DFFT_306_state_obs3(net1267_c1,net1267);
INTERCONNECT SplitCLK_6_345_SplitCLK_6_340(net1268_c1,net1268);
INTERCONNECT SplitCLK_6_345_SplitCLK_4_344(net1269_c1,net1269);
INTERCONNECT SplitCLK_4_344_SplitCLK_0_342(net1270_c1,net1270);
INTERCONNECT SplitCLK_4_344_SplitCLK_6_343(net1271_c1,net1271);
INTERCONNECT SplitCLK_6_343_SplitCLK_2_794(net1272_c1,net1272);
INTERCONNECT SplitCLK_6_343_SplitCLK_2_801(net1273_c1,net1273);
INTERCONNECT SplitCLK_0_342_SplitCLK_4_779(net1274_c1,net1274);
INTERCONNECT SplitCLK_0_342_SplitCLK_4_341(net1275_c1,net1275);
INTERCONNECT SplitCLK_4_341_AND2T_12_n36(net1276_c1,net1276);
INTERCONNECT SplitCLK_4_341_NOTT_120_n144(net1277_c1,net1277);
INTERCONNECT SplitCLK_6_340_SplitCLK_4_338(net1278_c1,net1278);
INTERCONNECT SplitCLK_6_340_SplitCLK_6_339(net1279_c1,net1279);
INTERCONNECT SplitCLK_6_339_SplitCLK_4_719(net1280_c1,net1280);
INTERCONNECT SplitCLK_6_339_SplitCLK_2_727(net1281_c1,net1281);
INTERCONNECT SplitCLK_4_338_SplitCLK_4_806(net1282_c1,net1282);
INTERCONNECT SplitCLK_4_338_SplitCLK_4_337(net1283_c1,net1283);
INTERCONNECT SplitCLK_4_337_DFFT_302__FPB_n758(net1284_c1,net1284);
INTERCONNECT SplitCLK_4_337_DFFT_303__FPB_n759(net1285_c1,net1285);
INTERCONNECT SplitCLK_0_336_SplitCLK_6_317(net1286_c1,net1286);
INTERCONNECT SplitCLK_0_336_SplitCLK_4_335(net1287_c1,net1287);
INTERCONNECT SplitCLK_4_335_SplitCLK_4_326(net1288_c1,net1288);
INTERCONNECT SplitCLK_4_335_SplitCLK_2_334(net1289_c1,net1289);
INTERCONNECT SplitCLK_2_334_SplitCLK_6_330(net1290_c1,net1290);
INTERCONNECT SplitCLK_2_334_SplitCLK_4_333(net1291_c1,net1291);
INTERCONNECT SplitCLK_4_333_SplitCLK_4_331(net1292_c1,net1292);
INTERCONNECT SplitCLK_4_333_SplitCLK_6_332(net1293_c1,net1293);
INTERCONNECT SplitCLK_6_332_SplitCLK_2_619(net1294_c1,net1294);
INTERCONNECT SplitCLK_6_332_SplitCLK_4_732(net1295_c1,net1295);
INTERCONNECT SplitCLK_4_331_SplitCLK_2_624(net1296_c1,net1296);
INTERCONNECT SplitCLK_4_331_SplitCLK_4_733(net1297_c1,net1297);
INTERCONNECT SplitCLK_6_330_SplitCLK_4_328(net1298_c1,net1298);
INTERCONNECT SplitCLK_6_330_SplitCLK_6_329(net1299_c1,net1299);
INTERCONNECT SplitCLK_6_329_SplitCLK_2_628(net1300_c1,net1300);
INTERCONNECT SplitCLK_6_329_SplitCLK_2_764(net1301_c1,net1301);
INTERCONNECT SplitCLK_4_328_SplitCLK_4_796(net1302_c1,net1302);
INTERCONNECT SplitCLK_4_328_SplitCLK_4_327(net1303_c1,net1303);
INTERCONNECT SplitCLK_4_327_NOTT_150_n198(net1304_c1,net1304);
INTERCONNECT SplitCLK_4_327_DFFT_169__FBL_n625(net1305_c1,net1305);
INTERCONNECT SplitCLK_4_326_SplitCLK_6_321(net1306_c1,net1306);
INTERCONNECT SplitCLK_4_326_SplitCLK_4_325(net1307_c1,net1307);
INTERCONNECT SplitCLK_4_325_SplitCLK_4_323(net1308_c1,net1308);
INTERCONNECT SplitCLK_4_325_SplitCLK_2_324(net1309_c1,net1309);
INTERCONNECT SplitCLK_2_324_SplitCLK_4_679(net1310_c1,net1310);
INTERCONNECT SplitCLK_2_324_SplitCLK_2_685(net1311_c1,net1311);
INTERCONNECT SplitCLK_4_323_SplitCLK_2_790(net1312_c1,net1312);
INTERCONNECT SplitCLK_4_323_SplitCLK_4_322(net1313_c1,net1313);
INTERCONNECT SplitCLK_4_322_DFFT_161__FBL_n617(net1314_c1,net1314);
INTERCONNECT SplitCLK_4_322_DFFT_249__FPB_n705(net1315_c1,net1315);
INTERCONNECT SplitCLK_6_321_SplitCLK_4_319(net1316_c1,net1316);
INTERCONNECT SplitCLK_6_321_SplitCLK_2_320(net1317_c1,net1317);
INTERCONNECT SplitCLK_2_320_SplitCLK_4_748(net1318_c1,net1318);
INTERCONNECT SplitCLK_2_320_SplitCLK_2_749(net1319_c1,net1319);
INTERCONNECT SplitCLK_4_319_SplitCLK_4_682(net1320_c1,net1320);
INTERCONNECT SplitCLK_4_319_SplitCLK_4_318(net1321_c1,net1321);
INTERCONNECT SplitCLK_4_318_AND2T_121_n145(net1322_c1,net1322);
INTERCONNECT SplitCLK_4_318_DFFT_172__FBL_n628(net1323_c1,net1323);
INTERCONNECT SplitCLK_6_317_SplitCLK_4_308(net1324_c1,net1324);
INTERCONNECT SplitCLK_6_317_SplitCLK_2_316(net1325_c1,net1325);
INTERCONNECT SplitCLK_2_316_SplitCLK_6_312(net1326_c1,net1326);
INTERCONNECT SplitCLK_2_316_SplitCLK_4_315(net1327_c1,net1327);
INTERCONNECT SplitCLK_4_315_SplitCLK_0_313(net1328_c1,net1328);
INTERCONNECT SplitCLK_4_315_SplitCLK_2_314(net1329_c1,net1329);
INTERCONNECT SplitCLK_2_314_SplitCLK_4_631(net1330_c1,net1330);
INTERCONNECT SplitCLK_2_314_SplitCLK_2_735(net1331_c1,net1331);
INTERCONNECT SplitCLK_0_313_SplitCLK_4_613(net1332_c1,net1332);
INTERCONNECT SplitCLK_0_313_SplitCLK_4_766(net1333_c1,net1333);
INTERCONNECT SplitCLK_6_312_SplitCLK_4_310(net1334_c1,net1334);
INTERCONNECT SplitCLK_6_312_SplitCLK_2_311(net1335_c1,net1335);
INTERCONNECT SplitCLK_2_311_SplitCLK_4_740(net1336_c1,net1336);
INTERCONNECT SplitCLK_2_311_SplitCLK_2_805(net1337_c1,net1337);
INTERCONNECT SplitCLK_4_310_SplitCLK_4_780(net1338_c1,net1338);
INTERCONNECT SplitCLK_4_310_SplitCLK_4_309(net1339_c1,net1339);
INTERCONNECT SplitCLK_4_309_AND2T_11_n35(net1340_c1,net1340);
INTERCONNECT SplitCLK_4_309_DFFT_157__PIPL_n211(net1341_c1,net1341);
INTERCONNECT SplitCLK_4_308_SplitCLK_6_303(net1342_c1,net1342);
INTERCONNECT SplitCLK_4_308_SplitCLK_6_307(net1343_c1,net1343);
INTERCONNECT SplitCLK_6_307_SplitCLK_0_305(net1344_c1,net1344);
INTERCONNECT SplitCLK_6_307_SplitCLK_2_306(net1345_c1,net1345);
INTERCONNECT SplitCLK_2_306_SplitCLK_2_745(net1346_c1,net1346);
INTERCONNECT SplitCLK_2_306_SplitCLK_4_768(net1347_c1,net1347);
INTERCONNECT SplitCLK_0_305_SplitCLK_4_772(net1348_c1,net1348);
INTERCONNECT SplitCLK_0_305_SplitCLK_4_304(net1349_c1,net1349);
INTERCONNECT SplitCLK_4_304_DFFT_253__FPB_n709(net1350_c1,net1350);
INTERCONNECT SplitCLK_4_304_DFFT_254__FPB_n710(net1351_c1,net1351);
INTERCONNECT SplitCLK_6_303_SplitCLK_4_301(net1352_c1,net1352);
INTERCONNECT SplitCLK_6_303_SplitCLK_6_302(net1353_c1,net1353);
INTERCONNECT SplitCLK_6_302_SplitCLK_4_714(net1354_c1,net1354);
INTERCONNECT SplitCLK_6_302_SplitCLK_2_787(net1355_c1,net1355);
INTERCONNECT SplitCLK_4_301_SplitCLK_4_759(net1356_c1,net1356);
INTERCONNECT SplitCLK_4_301_SplitCLK_4_300(net1357_c1,net1357);
INTERCONNECT SplitCLK_4_300_DFFT_300__FPB_n756(net1358_c1,net1358);
INTERCONNECT SplitCLK_4_300_DFFT_301__FPB_n757(net1359_c1,net1359);
INTERCONNECT GCLK_Pad_SplitCLK_0_810(GCLK_Pad,net1360);
INTERCONNECT Split_HOLD_943_NOTT_150_n198(net1361_c1,net1361);
INTERCONNECT Split_HOLD_944_DFFT_279__FPB_n735(net1362_c1,net1362);
INTERCONNECT Split_HOLD_945_XOR2T_45_n69(net1363_c1,net1363);

endmodule
