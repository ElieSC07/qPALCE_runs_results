module TAP_half_route(
input GCLK_Pad,
input TMS_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output output1_Pad);

wire net0_c1;
wire state_obs0_Pad;
wire net1_c1;
wire state_obs1_Pad;
wire TMS_Pad;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire TRST_Pad;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire output1_Pad;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire GCLK_Pad;
wire net184;

NOTT NOTT_7_n22(net109,net64,net4_c1);
NOTT NOTT_8_n23(net182,net55,net6_c1);
NOTT NOTT_9_n24(net108,net62,net9_c1);
AND2T AND2T_10_n25(net107,net50,net48,net12_c1);
AND2T AND2T_21_n36(net106,net29,net35,net20_c1);
AND2T AND2T_30_n45(net164,net19,net79,net22_c1);
AND2T AND2T_22_n37(net105,net58,net17,net23_c1);
AND2T AND2T_14_n29(net126,net21,net54,net24_c1);
AND2T AND2T_23_n38(net104,net23,net14,net26_c1);
AND2T AND2T_16_n31(net103,net57,net72,net5_c1);
AND2T AND2T_25_n40(net174,net38,net75,net7_c1);
AND2T AND2T_17_n32(net102,net5,net52,net8_c1);
AND2T AND2T_26_n41(net144,net7,net33,net10_c1);
AND2T AND2T_18_n33(net136,net60,net31,net11_c1);
AND2T AND2T_27_n42(net101,net39,net76,net13_c1);
AND2T AND2T_28_n43(net100,net4,net77,net16_c1);
DFFT DFFT_32__FBL_n74(net156,net8,net66_c1);
DFFT DFFT_40__FPB_n82(net99,net80,net73_c1);
DFFT DFFT_33__FBL_n75(net137,net26,net67_c1);
DFFT DFFT_41__FPB_n83(net98,net73,net74_c1);
DFFT DFFT_34__FBL_n76(net97,net10,net68_c1);
DFFT DFFT_42__FPB_n84(net175,net27,net75_c1);
DFFT DFFT_35__FBL_n77(net96,net78,net69_c1);
DFFT DFFT_43__FPB_n85(net95,net42,net76_c1);
OR2T OR2T_11_n26(net94,net51,net71,net15_c1);
OR2T OR2T_20_n35(net93,net41,net49,net17_c1);
DFFT DFFT_36__FBL_n78(net92,net22,net70_c1);
OR2T OR2T_13_n28(net91,net45,net43,net21_c1);
OR2T OR2T_15_n30(net90,net65,net37,net3_c1);
OR2T OR2T_24_n39(net89,net81,net47,net27_c1);
OR2T OR2T_19_n34(net145,net11,net74,net14_c1);
OR2T OR2T_29_n44(net157,net16,net32,net19_c1);
DFFT DFFT_44__FPB_n86(net183,net28,net77_c1);
DFFT DFFT_45__FPB_n87(net165,net56,net79_c1);
DFFT DFFT_37__FPB_n79(net88,net13,net78_c1);
DFFT DFFT_38__FPB_n80(net87,net61,net71_c1);
DFFT DFFT_39__FPB_n81(net86,net3,net72_c1);
NOTT NOTT_12_n27(net85,net46,net18_c1);
NOTT NOTT_31_n46(net127,net63,net25_c1);
SPLITT Split_62_state_obs0(net67,net80_c1,net0_c1);
SPLITT Split_63_state_obs1(net68,net81_c1,net1_c1);
SPLITT Split_61_output1(net66,net65_c1,net82_c1);
SPLITT Split_60_n102(net40,net42_c1,net61_c1);
SPLITT Split_64_n106(net69,net43_c1,net62_c1);
SPLITT Split_65_n107(net70,net44_c1,net63_c1);
SPLITT Split_58_n100(net25,net40_c1,net59_c1);
SPLITT Split_66_n108(net44,net45_c1,net64_c1);
SPLITT Split_59_n101(net59,net41_c1,net60_c1);
SPLITT Split_50_n92(net9,net30_c1,net49_c1);
SPLITT Split_51_n93(net30,net31_c1,net50_c1);
SPLITT Split_52_n94(net12,net32_c1,net51_c1);
SPLITT Split_53_n95(net15,net33_c1,net52_c1);
SPLITT Split_46_n88(net2,net34_c1,net53_c1);
SPLITT Split_54_n96(net18,net35_c1,net54_c1);
SPLITT Split_47_n89(net53,net37_c1,net55_c1);
SPLITT Split_55_n97(net24,net36_c1,net56_c1);
SPLITT Split_48_n90(net34,net28_c1,net47_c1);
SPLITT Split_56_n98(net36,net38_c1,net57_c1);
SPLITT Split_49_n91(net6,net29_c1,net48_c1);
SPLITT Split_57_n99(net20,net39_c1,net58_c1);
SPLITT SplitCLK_4_40(net181,net182_c1,net183_c1);
SPLITT SplitCLK_6_41(net176,net181_c1,net180_c1);
SPLITT SplitCLK_0_42(net177,net178_c1,net179_c1);
SPLITT SplitCLK_4_43(net166,net176_c1,net177_c1);
SPLITT SplitCLK_4_44(net173,net174_c1,net175_c1);
SPLITT SplitCLK_6_45(net168,net173_c1,net172_c1);
SPLITT SplitCLK_6_46(net169,net170_c1,net171_c1);
SPLITT SplitCLK_6_47(net167,net168_c1,net169_c1);
SPLITT SplitCLK_6_48(net146,net166_c1,net167_c1);
SPLITT SplitCLK_4_49(net163,net164_c1,net165_c1);
SPLITT SplitCLK_0_50(net158,net162_c1,net163_c1);
SPLITT SplitCLK_4_51(net159,net160_c1,net161_c1);
SPLITT SplitCLK_4_52(net148,net158_c1,net159_c1);
SPLITT SplitCLK_4_53(net155,net156_c1,net157_c1);
SPLITT SplitCLK_0_54(net150,net154_c1,net155_c1);
SPLITT SplitCLK_4_55(net151,net152_c1,net153_c1);
SPLITT SplitCLK_6_56(net149,net150_c1,net151_c1);
SPLITT SplitCLK_4_57(net147,net149_c1,net148_c1);
SPLITT SplitCLK_0_58(net83,net146_c1,net147_c1);
SPLITT SplitCLK_4_59(net143,net145_c1,net144_c1);
SPLITT SplitCLK_0_60(net138,net142_c1,net143_c1);
SPLITT SplitCLK_2_61(net139,net141_c1,net140_c1);
SPLITT SplitCLK_4_62(net128,net139_c1,net138_c1);
SPLITT SplitCLK_4_63(net135,net136_c1,net137_c1);
SPLITT SplitCLK_2_64(net130,net134_c1,net135_c1);
SPLITT SplitCLK_2_65(net131,net132_c1,net133_c1);
SPLITT SplitCLK_6_66(net129,net130_c1,net131_c1);
SPLITT SplitCLK_6_67(net110,net128_c1,net129_c1);
SPLITT SplitCLK_4_68(net125,net127_c1,net126_c1);
SPLITT SplitCLK_6_69(net120,net125_c1,net124_c1);
SPLITT SplitCLK_0_70(net121,net123_c1,net122_c1);
SPLITT SplitCLK_4_71(net112,net120_c1,net121_c1);
SPLITT SplitCLK_0_72(net114,net118_c1,net119_c1);
SPLITT SplitCLK_0_73(net115,net116_c1,net117_c1);
SPLITT SplitCLK_2_74(net113,net115_c1,net114_c1);
SPLITT SplitCLK_4_75(net111,net113_c1,net112_c1);
SPLITT SplitCLK_2_76(net84,net111_c1,net110_c1);
wire dummy0;
SPLITT SplitCLK_2_77(net162,net109_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_4_78(net132,net108_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_79(net178,net107_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_4_80(net170,net106_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_81(net133,net105_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_2_82(net142,net104_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_4_83(net122,net103_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_2_84(net152,net102_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_2_85(net118,net101_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_4_86(net179,net100_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_2_87(net134,net99_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_2_88(net172,net98_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_2_89(net140,net97_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_4_90(net119,net96_c1,dummy13);
wire dummy14;
SPLITT SplitCLK_2_91(net124,net95_c1,dummy14);
wire dummy15;
SPLITT SplitCLK_2_92(net154,net94_c1,dummy15);
wire dummy16;
SPLITT SplitCLK_4_93(net141,net93_c1,dummy16);
wire dummy17;
SPLITT SplitCLK_2_94(net160,net92_c1,dummy17);
wire dummy18;
SPLITT SplitCLK_2_95(net123,net91_c1,dummy18);
wire dummy19;
SPLITT SplitCLK_4_96(net161,net90_c1,dummy19);
wire dummy20;
SPLITT SplitCLK_2_97(net180,net89_c1,dummy20);
wire dummy21;
SPLITT SplitCLK_2_98(net116,net88_c1,dummy21);
wire dummy22;
SPLITT SplitCLK_4_99(net171,net87_c1,dummy22);
wire dummy23;
SPLITT SplitCLK_4_100(net153,net86_c1,dummy23);
wire dummy24;
SPLITT SplitCLK_4_101(net117,net85_c1,dummy24);
SPLITT SplitCLK_0_102(net184,net83_c1,net84_c1);
INTERCONNECT Split_62_state_obs0_state_obs0_Pad(net0_c1,state_obs0_Pad);
INTERCONNECT Split_63_state_obs1_state_obs1_Pad(net1_c1,state_obs1_Pad);
INTERCONNECT TMS_Pad_Split_46_n88(TMS_Pad,net2);
INTERCONNECT OR2T_15_n30_DFFT_39__FPB_n81(net3_c1,net3);
INTERCONNECT NOTT_7_n22_AND2T_28_n43(net4_c1,net4);
INTERCONNECT AND2T_16_n31_AND2T_17_n32(net5_c1,net5);
INTERCONNECT NOTT_8_n23_Split_49_n91(net6_c1,net6);
INTERCONNECT AND2T_25_n40_AND2T_26_n41(net7_c1,net7);
INTERCONNECT AND2T_17_n32_DFFT_32__FBL_n74(net8_c1,net8);
INTERCONNECT NOTT_9_n24_Split_50_n92(net9_c1,net9);
INTERCONNECT AND2T_26_n41_DFFT_34__FBL_n76(net10_c1,net10);
INTERCONNECT AND2T_18_n33_OR2T_19_n34(net11_c1,net11);
INTERCONNECT AND2T_10_n25_Split_52_n94(net12_c1,net12);
INTERCONNECT AND2T_27_n42_DFFT_37__FPB_n79(net13_c1,net13);
INTERCONNECT OR2T_19_n34_AND2T_23_n38(net14_c1,net14);
INTERCONNECT OR2T_11_n26_Split_53_n95(net15_c1,net15);
INTERCONNECT AND2T_28_n43_OR2T_29_n44(net16_c1,net16);
INTERCONNECT OR2T_20_n35_AND2T_22_n37(net17_c1,net17);
INTERCONNECT NOTT_12_n27_Split_54_n96(net18_c1,net18);
INTERCONNECT OR2T_29_n44_AND2T_30_n45(net19_c1,net19);
INTERCONNECT AND2T_21_n36_Split_57_n99(net20_c1,net20);
INTERCONNECT OR2T_13_n28_AND2T_14_n29(net21_c1,net21);
INTERCONNECT AND2T_30_n45_DFFT_36__FBL_n78(net22_c1,net22);
INTERCONNECT AND2T_22_n37_AND2T_23_n38(net23_c1,net23);
INTERCONNECT AND2T_14_n29_Split_55_n97(net24_c1,net24);
INTERCONNECT NOTT_31_n46_Split_58_n100(net25_c1,net25);
INTERCONNECT AND2T_23_n38_DFFT_33__FBL_n75(net26_c1,net26);
INTERCONNECT OR2T_24_n39_DFFT_42__FPB_n84(net27_c1,net27);
INTERCONNECT Split_48_n90_DFFT_44__FPB_n86(net28_c1,net28);
INTERCONNECT Split_49_n91_AND2T_21_n36(net29_c1,net29);
INTERCONNECT Split_50_n92_Split_51_n93(net30_c1,net30);
INTERCONNECT Split_51_n93_AND2T_18_n33(net31_c1,net31);
INTERCONNECT Split_52_n94_OR2T_29_n44(net32_c1,net32);
INTERCONNECT Split_53_n95_AND2T_26_n41(net33_c1,net33);
INTERCONNECT Split_46_n88_Split_48_n90(net34_c1,net34);
INTERCONNECT Split_54_n96_AND2T_21_n36(net35_c1,net35);
INTERCONNECT Split_55_n97_Split_56_n98(net36_c1,net36);
INTERCONNECT Split_47_n89_OR2T_15_n30(net37_c1,net37);
INTERCONNECT Split_56_n98_AND2T_25_n40(net38_c1,net38);
INTERCONNECT Split_57_n99_AND2T_27_n42(net39_c1,net39);
INTERCONNECT Split_58_n100_Split_60_n102(net40_c1,net40);
INTERCONNECT Split_59_n101_OR2T_20_n35(net41_c1,net41);
INTERCONNECT Split_60_n102_DFFT_43__FPB_n85(net42_c1,net42);
INTERCONNECT Split_64_n106_OR2T_13_n28(net43_c1,net43);
INTERCONNECT Split_65_n107_Split_66_n108(net44_c1,net44);
INTERCONNECT Split_66_n108_OR2T_13_n28(net45_c1,net45);
INTERCONNECT TRST_Pad_NOTT_12_n27(TRST_Pad,net46);
INTERCONNECT Split_48_n90_OR2T_24_n39(net47_c1,net47);
INTERCONNECT Split_49_n91_AND2T_10_n25(net48_c1,net48);
INTERCONNECT Split_50_n92_OR2T_20_n35(net49_c1,net49);
INTERCONNECT Split_51_n93_AND2T_10_n25(net50_c1,net50);
INTERCONNECT Split_52_n94_OR2T_11_n26(net51_c1,net51);
INTERCONNECT Split_53_n95_AND2T_17_n32(net52_c1,net52);
INTERCONNECT Split_46_n88_Split_47_n89(net53_c1,net53);
INTERCONNECT Split_54_n96_AND2T_14_n29(net54_c1,net54);
INTERCONNECT Split_47_n89_NOTT_8_n23(net55_c1,net55);
INTERCONNECT Split_55_n97_DFFT_45__FPB_n87(net56_c1,net56);
INTERCONNECT Split_56_n98_AND2T_16_n31(net57_c1,net57);
INTERCONNECT Split_57_n99_AND2T_22_n37(net58_c1,net58);
INTERCONNECT Split_58_n100_Split_59_n101(net59_c1,net59);
INTERCONNECT Split_59_n101_AND2T_18_n33(net60_c1,net60);
INTERCONNECT Split_60_n102_DFFT_38__FPB_n80(net61_c1,net61);
INTERCONNECT Split_64_n106_NOTT_9_n24(net62_c1,net62);
INTERCONNECT Split_65_n107_NOTT_31_n46(net63_c1,net63);
INTERCONNECT Split_66_n108_NOTT_7_n22(net64_c1,net64);
INTERCONNECT Split_61_output1_OR2T_15_n30(net65_c1,net65);
INTERCONNECT DFFT_32__FBL_n74_Split_61_output1(net66_c1,net66);
INTERCONNECT DFFT_33__FBL_n75_Split_62_state_obs0(net67_c1,net67);
INTERCONNECT DFFT_34__FBL_n76_Split_63_state_obs1(net68_c1,net68);
INTERCONNECT DFFT_35__FBL_n77_Split_64_n106(net69_c1,net69);
INTERCONNECT DFFT_36__FBL_n78_Split_65_n107(net70_c1,net70);
INTERCONNECT DFFT_38__FPB_n80_OR2T_11_n26(net71_c1,net71);
INTERCONNECT DFFT_39__FPB_n81_AND2T_16_n31(net72_c1,net72);
INTERCONNECT DFFT_40__FPB_n82_DFFT_41__FPB_n83(net73_c1,net73);
INTERCONNECT DFFT_41__FPB_n83_OR2T_19_n34(net74_c1,net74);
INTERCONNECT DFFT_42__FPB_n84_AND2T_25_n40(net75_c1,net75);
INTERCONNECT DFFT_43__FPB_n85_AND2T_27_n42(net76_c1,net76);
INTERCONNECT DFFT_44__FPB_n86_AND2T_28_n43(net77_c1,net77);
INTERCONNECT DFFT_37__FPB_n79_DFFT_35__FBL_n77(net78_c1,net78);
INTERCONNECT DFFT_45__FPB_n87_AND2T_30_n45(net79_c1,net79);
INTERCONNECT Split_62_state_obs0_DFFT_40__FPB_n82(net80_c1,net80);
INTERCONNECT Split_63_state_obs1_OR2T_24_n39(net81_c1,net81);
INTERCONNECT Split_61_output1_output1_Pad(net82_c1,output1_Pad);
INTERCONNECT SplitCLK_0_102_SplitCLK_0_58(net83_c1,net83);
INTERCONNECT SplitCLK_0_102_SplitCLK_2_76(net84_c1,net84);
INTERCONNECT SplitCLK_4_101_NOTT_12_n27(net85_c1,net85);
INTERCONNECT SplitCLK_4_100_DFFT_39__FPB_n81(net86_c1,net86);
INTERCONNECT SplitCLK_4_99_DFFT_38__FPB_n80(net87_c1,net87);
INTERCONNECT SplitCLK_2_98_DFFT_37__FPB_n79(net88_c1,net88);
INTERCONNECT SplitCLK_2_97_OR2T_24_n39(net89_c1,net89);
INTERCONNECT SplitCLK_4_96_OR2T_15_n30(net90_c1,net90);
INTERCONNECT SplitCLK_2_95_OR2T_13_n28(net91_c1,net91);
INTERCONNECT SplitCLK_2_94_DFFT_36__FBL_n78(net92_c1,net92);
INTERCONNECT SplitCLK_4_93_OR2T_20_n35(net93_c1,net93);
INTERCONNECT SplitCLK_2_92_OR2T_11_n26(net94_c1,net94);
INTERCONNECT SplitCLK_2_91_DFFT_43__FPB_n85(net95_c1,net95);
INTERCONNECT SplitCLK_4_90_DFFT_35__FBL_n77(net96_c1,net96);
INTERCONNECT SplitCLK_2_89_DFFT_34__FBL_n76(net97_c1,net97);
INTERCONNECT SplitCLK_2_88_DFFT_41__FPB_n83(net98_c1,net98);
INTERCONNECT SplitCLK_2_87_DFFT_40__FPB_n82(net99_c1,net99);
INTERCONNECT SplitCLK_4_86_AND2T_28_n43(net100_c1,net100);
INTERCONNECT SplitCLK_2_85_AND2T_27_n42(net101_c1,net101);
INTERCONNECT SplitCLK_2_84_AND2T_17_n32(net102_c1,net102);
INTERCONNECT SplitCLK_4_83_AND2T_16_n31(net103_c1,net103);
INTERCONNECT SplitCLK_2_82_AND2T_23_n38(net104_c1,net104);
INTERCONNECT SplitCLK_2_81_AND2T_22_n37(net105_c1,net105);
INTERCONNECT SplitCLK_4_80_AND2T_21_n36(net106_c1,net106);
INTERCONNECT SplitCLK_2_79_AND2T_10_n25(net107_c1,net107);
INTERCONNECT SplitCLK_4_78_NOTT_9_n24(net108_c1,net108);
INTERCONNECT SplitCLK_2_77_NOTT_7_n22(net109_c1,net109);
INTERCONNECT SplitCLK_2_76_SplitCLK_6_67(net110_c1,net110);
INTERCONNECT SplitCLK_2_76_SplitCLK_4_75(net111_c1,net111);
INTERCONNECT SplitCLK_4_75_SplitCLK_4_71(net112_c1,net112);
INTERCONNECT SplitCLK_4_75_SplitCLK_2_74(net113_c1,net113);
INTERCONNECT SplitCLK_2_74_SplitCLK_0_72(net114_c1,net114);
INTERCONNECT SplitCLK_2_74_SplitCLK_0_73(net115_c1,net115);
INTERCONNECT SplitCLK_0_73_SplitCLK_2_98(net116_c1,net116);
INTERCONNECT SplitCLK_0_73_SplitCLK_4_101(net117_c1,net117);
INTERCONNECT SplitCLK_0_72_SplitCLK_2_85(net118_c1,net118);
INTERCONNECT SplitCLK_0_72_SplitCLK_4_90(net119_c1,net119);
INTERCONNECT SplitCLK_4_71_SplitCLK_6_69(net120_c1,net120);
INTERCONNECT SplitCLK_4_71_SplitCLK_0_70(net121_c1,net121);
INTERCONNECT SplitCLK_0_70_SplitCLK_4_83(net122_c1,net122);
INTERCONNECT SplitCLK_0_70_SplitCLK_2_95(net123_c1,net123);
INTERCONNECT SplitCLK_6_69_SplitCLK_2_91(net124_c1,net124);
INTERCONNECT SplitCLK_6_69_SplitCLK_4_68(net125_c1,net125);
INTERCONNECT SplitCLK_4_68_AND2T_14_n29(net126_c1,net126);
INTERCONNECT SplitCLK_4_68_NOTT_31_n46(net127_c1,net127);
INTERCONNECT SplitCLK_6_67_SplitCLK_4_62(net128_c1,net128);
INTERCONNECT SplitCLK_6_67_SplitCLK_6_66(net129_c1,net129);
INTERCONNECT SplitCLK_6_66_SplitCLK_2_64(net130_c1,net130);
INTERCONNECT SplitCLK_6_66_SplitCLK_2_65(net131_c1,net131);
INTERCONNECT SplitCLK_2_65_SplitCLK_4_78(net132_c1,net132);
INTERCONNECT SplitCLK_2_65_SplitCLK_2_81(net133_c1,net133);
INTERCONNECT SplitCLK_2_64_SplitCLK_2_87(net134_c1,net134);
INTERCONNECT SplitCLK_2_64_SplitCLK_4_63(net135_c1,net135);
INTERCONNECT SplitCLK_4_63_AND2T_18_n33(net136_c1,net136);
INTERCONNECT SplitCLK_4_63_DFFT_33__FBL_n75(net137_c1,net137);
INTERCONNECT SplitCLK_4_62_SplitCLK_0_60(net138_c1,net138);
INTERCONNECT SplitCLK_4_62_SplitCLK_2_61(net139_c1,net139);
INTERCONNECT SplitCLK_2_61_SplitCLK_2_89(net140_c1,net140);
INTERCONNECT SplitCLK_2_61_SplitCLK_4_93(net141_c1,net141);
INTERCONNECT SplitCLK_0_60_SplitCLK_2_82(net142_c1,net142);
INTERCONNECT SplitCLK_0_60_SplitCLK_4_59(net143_c1,net143);
INTERCONNECT SplitCLK_4_59_AND2T_26_n41(net144_c1,net144);
INTERCONNECT SplitCLK_4_59_OR2T_19_n34(net145_c1,net145);
INTERCONNECT SplitCLK_0_58_SplitCLK_6_48(net146_c1,net146);
INTERCONNECT SplitCLK_0_58_SplitCLK_4_57(net147_c1,net147);
INTERCONNECT SplitCLK_4_57_SplitCLK_4_52(net148_c1,net148);
INTERCONNECT SplitCLK_4_57_SplitCLK_6_56(net149_c1,net149);
INTERCONNECT SplitCLK_6_56_SplitCLK_0_54(net150_c1,net150);
INTERCONNECT SplitCLK_6_56_SplitCLK_4_55(net151_c1,net151);
INTERCONNECT SplitCLK_4_55_SplitCLK_2_84(net152_c1,net152);
INTERCONNECT SplitCLK_4_55_SplitCLK_4_100(net153_c1,net153);
INTERCONNECT SplitCLK_0_54_SplitCLK_2_92(net154_c1,net154);
INTERCONNECT SplitCLK_0_54_SplitCLK_4_53(net155_c1,net155);
INTERCONNECT SplitCLK_4_53_DFFT_32__FBL_n74(net156_c1,net156);
INTERCONNECT SplitCLK_4_53_OR2T_29_n44(net157_c1,net157);
INTERCONNECT SplitCLK_4_52_SplitCLK_0_50(net158_c1,net158);
INTERCONNECT SplitCLK_4_52_SplitCLK_4_51(net159_c1,net159);
INTERCONNECT SplitCLK_4_51_SplitCLK_2_94(net160_c1,net160);
INTERCONNECT SplitCLK_4_51_SplitCLK_4_96(net161_c1,net161);
INTERCONNECT SplitCLK_0_50_SplitCLK_2_77(net162_c1,net162);
INTERCONNECT SplitCLK_0_50_SplitCLK_4_49(net163_c1,net163);
INTERCONNECT SplitCLK_4_49_AND2T_30_n45(net164_c1,net164);
INTERCONNECT SplitCLK_4_49_DFFT_45__FPB_n87(net165_c1,net165);
INTERCONNECT SplitCLK_6_48_SplitCLK_4_43(net166_c1,net166);
INTERCONNECT SplitCLK_6_48_SplitCLK_6_47(net167_c1,net167);
INTERCONNECT SplitCLK_6_47_SplitCLK_6_45(net168_c1,net168);
INTERCONNECT SplitCLK_6_47_SplitCLK_6_46(net169_c1,net169);
INTERCONNECT SplitCLK_6_46_SplitCLK_4_80(net170_c1,net170);
INTERCONNECT SplitCLK_6_46_SplitCLK_4_99(net171_c1,net171);
INTERCONNECT SplitCLK_6_45_SplitCLK_2_88(net172_c1,net172);
INTERCONNECT SplitCLK_6_45_SplitCLK_4_44(net173_c1,net173);
INTERCONNECT SplitCLK_4_44_AND2T_25_n40(net174_c1,net174);
INTERCONNECT SplitCLK_4_44_DFFT_42__FPB_n84(net175_c1,net175);
INTERCONNECT SplitCLK_4_43_SplitCLK_6_41(net176_c1,net176);
INTERCONNECT SplitCLK_4_43_SplitCLK_0_42(net177_c1,net177);
INTERCONNECT SplitCLK_0_42_SplitCLK_2_79(net178_c1,net178);
INTERCONNECT SplitCLK_0_42_SplitCLK_4_86(net179_c1,net179);
INTERCONNECT SplitCLK_6_41_SplitCLK_2_97(net180_c1,net180);
INTERCONNECT SplitCLK_6_41_SplitCLK_4_40(net181_c1,net181);
INTERCONNECT SplitCLK_4_40_NOTT_8_n23(net182_c1,net182);
INTERCONNECT SplitCLK_4_40_DFFT_44__FPB_n86(net183_c1,net183);
INTERCONNECT GCLK_Pad_SplitCLK_0_102(GCLK_Pad,net184);

endmodule
