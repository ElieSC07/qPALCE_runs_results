module KSA2_route(
input GCLK_Pad,
input a0_Pad,
input a1_Pad,
input b0_Pad,
input b1_Pad,
input cin_Pad,
output cout_Pad,
output sum0_Pad,
output sum1_Pad);

wire a0_Pad;
wire net0;
wire a1_Pad;
wire net1;
wire b0_Pad;
wire net2;
wire b1_Pad;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire cin_Pad;
wire net24;
wire net25_c1;
wire cout_Pad;
wire net26_c1;
wire sum0_Pad;
wire net27_c1;
wire sum1_Pad;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire GCLK_Pad;
wire net97;

XOR2T XOR2T_10_n10(net85,net30,net44,net5_c1);
XOR2T XOR2T_11_n11(net75,net28,net36,net6_c1);
XOR2T XOR2T_15_sum1(net86,net9,net40,net27_c1);
XOR2T XOR2T_9_n9(net95,net37,net34,net4_c1);
AND2T AND2T_12_n12(net58,net16,net45,net7_c1);
AND2T AND2T_13_n13(net91,net23,net20,net8_c1);
AND2T AND2T_16_n16(net57,net19,net41,net10_c1);
AND2T AND2T_17_n17(net92,net35,net32,net11_c1);
AND2T AND2T_18_n18(net56,net14,net22,net12_c1);
DFFT DFFT_21__FPB_n48(net55,net29,net44_c1);
DFFT DFFT_22__FPB_n49(net96,net15,net45_c1);
DFFT DFFT_23__FPB_n50(net54,net21,net38_c1);
DFFT DFFT_24__FPB_n51(net67,net18,net39_c1);
DFFT DFFT_25__FPB_n52(net53,net39,net40_c1);
DFFT DFFT_26__FPB_n53(net76,net31,net41_c1);
DFFT DFFT_27__FPB_n54(net52,net12,net42_c1);
OR2T OR2T_14_n14(net51,net33,net38,net9_c1);
OR2T OR2T_19_n19(net50,net11,net42,net13_c1);
DFFT DFFT_28__FPB_n55(net68,net5,net43_c1);
DFFT DFFT_29_sum0(net49,net43,net26_c1);
OR2T OR2T_20_cout(net48,net13,net10,net25_c1);
SPLITT Split_30_n57(net0,net20_c1,net34_c1);
SPLITT Split_31_n58(net1,net22_c1,net36_c1);
SPLITT Split_32_n59(net2,net23_c1,net37_c1);
SPLITT Split_33_n60(net3,net14_c1,net28_c1);
SPLITT Split_34_n61(net24,net15_c1,net29_c1);
SPLITT Split_35_n62(net4,net16_c1,net30_c1);
SPLITT Split_36_n63(net6,net17_c1,net31_c1);
SPLITT Split_37_n64(net17,net18_c1,net32_c1);
SPLITT Split_38_n65(net7,net19_c1,net33_c1);
SPLITT Split_39_n66(net8,net21_c1,net35_c1);
SPLITT SplitCLK_4_22(net94,net95_c1,net96_c1);
SPLITT SplitCLK_4_23(net87,net94_c1,net93_c1);
SPLITT SplitCLK_4_24(net90,net91_c1,net92_c1);
SPLITT SplitCLK_2_25(net88,net89_c1,net90_c1);
SPLITT SplitCLK_6_26(net77,net87_c1,net88_c1);
SPLITT SplitCLK_4_27(net84,net86_c1,net85_c1);
SPLITT SplitCLK_4_28(net79,net83_c1,net84_c1);
SPLITT SplitCLK_2_29(net80,net82_c1,net81_c1);
SPLITT SplitCLK_4_30(net78,net80_c1,net79_c1);
SPLITT SplitCLK_0_31(net46,net77_c1,net78_c1);
SPLITT SplitCLK_4_32(net74,net75_c1,net76_c1);
SPLITT SplitCLK_4_33(net69,net73_c1,net74_c1);
SPLITT SplitCLK_6_34(net70,net71_c1,net72_c1);
SPLITT SplitCLK_6_35(net59,net69_c1,net70_c1);
SPLITT SplitCLK_4_36(net66,net67_c1,net68_c1);
SPLITT SplitCLK_2_37(net61,net65_c1,net66_c1);
SPLITT SplitCLK_6_38(net62,net63_c1,net64_c1);
SPLITT SplitCLK_4_39(net60,net62_c1,net61_c1);
SPLITT SplitCLK_2_40(net47,net60_c1,net59_c1);
wire dummy0;
SPLITT SplitCLK_4_41(net89,net58_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_2_42(net63,net57_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_43(net71,net56_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_4_44(net93,net55_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_45(net81,net54_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_4_46(net82,net53_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_4_47(net72,net52_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_2_48(net83,net51_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_2_49(net73,net50_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_4_50(net64,net49_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_2_51(net65,net48_c1,dummy10);
SPLITT SplitCLK_0_52(net97,net46_c1,net47_c1);
INTERCONNECT a0_Pad_Split_30_n57(a0_Pad,net0);
INTERCONNECT a1_Pad_Split_31_n58(a1_Pad,net1);
INTERCONNECT b0_Pad_Split_32_n59(b0_Pad,net2);
INTERCONNECT b1_Pad_Split_33_n60(b1_Pad,net3);
INTERCONNECT XOR2T_9_n9_Split_35_n62(net4_c1,net4);
INTERCONNECT XOR2T_10_n10_DFFT_28__FPB_n55(net5_c1,net5);
INTERCONNECT XOR2T_11_n11_Split_36_n63(net6_c1,net6);
INTERCONNECT AND2T_12_n12_Split_38_n65(net7_c1,net7);
INTERCONNECT AND2T_13_n13_Split_39_n66(net8_c1,net8);
INTERCONNECT OR2T_14_n14_XOR2T_15_sum1(net9_c1,net9);
INTERCONNECT AND2T_16_n16_OR2T_20_cout(net10_c1,net10);
INTERCONNECT AND2T_17_n17_OR2T_19_n19(net11_c1,net11);
INTERCONNECT AND2T_18_n18_DFFT_27__FPB_n54(net12_c1,net12);
INTERCONNECT OR2T_19_n19_OR2T_20_cout(net13_c1,net13);
INTERCONNECT Split_33_n60_AND2T_18_n18(net14_c1,net14);
INTERCONNECT Split_34_n61_DFFT_22__FPB_n49(net15_c1,net15);
INTERCONNECT Split_35_n62_AND2T_12_n12(net16_c1,net16);
INTERCONNECT Split_36_n63_Split_37_n64(net17_c1,net17);
INTERCONNECT Split_37_n64_DFFT_24__FPB_n51(net18_c1,net18);
INTERCONNECT Split_38_n65_AND2T_16_n16(net19_c1,net19);
INTERCONNECT Split_30_n57_AND2T_13_n13(net20_c1,net20);
INTERCONNECT Split_39_n66_DFFT_23__FPB_n50(net21_c1,net21);
INTERCONNECT Split_31_n58_AND2T_18_n18(net22_c1,net22);
INTERCONNECT Split_32_n59_AND2T_13_n13(net23_c1,net23);
INTERCONNECT cin_Pad_Split_34_n61(cin_Pad,net24);
INTERCONNECT OR2T_20_cout_cout_Pad(net25_c1,cout_Pad);
INTERCONNECT DFFT_29_sum0_sum0_Pad(net26_c1,sum0_Pad);
INTERCONNECT XOR2T_15_sum1_sum1_Pad(net27_c1,sum1_Pad);
INTERCONNECT Split_33_n60_XOR2T_11_n11(net28_c1,net28);
INTERCONNECT Split_34_n61_DFFT_21__FPB_n48(net29_c1,net29);
INTERCONNECT Split_35_n62_XOR2T_10_n10(net30_c1,net30);
INTERCONNECT Split_36_n63_DFFT_26__FPB_n53(net31_c1,net31);
INTERCONNECT Split_37_n64_AND2T_17_n17(net32_c1,net32);
INTERCONNECT Split_38_n65_OR2T_14_n14(net33_c1,net33);
INTERCONNECT Split_30_n57_XOR2T_9_n9(net34_c1,net34);
INTERCONNECT Split_39_n66_AND2T_17_n17(net35_c1,net35);
INTERCONNECT Split_31_n58_XOR2T_11_n11(net36_c1,net36);
INTERCONNECT Split_32_n59_XOR2T_9_n9(net37_c1,net37);
INTERCONNECT DFFT_23__FPB_n50_OR2T_14_n14(net38_c1,net38);
INTERCONNECT DFFT_24__FPB_n51_DFFT_25__FPB_n52(net39_c1,net39);
INTERCONNECT DFFT_25__FPB_n52_XOR2T_15_sum1(net40_c1,net40);
INTERCONNECT DFFT_26__FPB_n53_AND2T_16_n16(net41_c1,net41);
INTERCONNECT DFFT_27__FPB_n54_OR2T_19_n19(net42_c1,net42);
INTERCONNECT DFFT_28__FPB_n55_DFFT_29_sum0(net43_c1,net43);
INTERCONNECT DFFT_21__FPB_n48_XOR2T_10_n10(net44_c1,net44);
INTERCONNECT DFFT_22__FPB_n49_AND2T_12_n12(net45_c1,net45);
INTERCONNECT SplitCLK_0_52_SplitCLK_0_31(net46_c1,net46);
INTERCONNECT SplitCLK_0_52_SplitCLK_2_40(net47_c1,net47);
INTERCONNECT SplitCLK_2_51_OR2T_20_cout(net48_c1,net48);
INTERCONNECT SplitCLK_4_50_DFFT_29_sum0(net49_c1,net49);
INTERCONNECT SplitCLK_2_49_OR2T_19_n19(net50_c1,net50);
INTERCONNECT SplitCLK_2_48_OR2T_14_n14(net51_c1,net51);
INTERCONNECT SplitCLK_4_47_DFFT_27__FPB_n54(net52_c1,net52);
INTERCONNECT SplitCLK_4_46_DFFT_25__FPB_n52(net53_c1,net53);
INTERCONNECT SplitCLK_2_45_DFFT_23__FPB_n50(net54_c1,net54);
INTERCONNECT SplitCLK_4_44_DFFT_21__FPB_n48(net55_c1,net55);
INTERCONNECT SplitCLK_2_43_AND2T_18_n18(net56_c1,net56);
INTERCONNECT SplitCLK_2_42_AND2T_16_n16(net57_c1,net57);
INTERCONNECT SplitCLK_4_41_AND2T_12_n12(net58_c1,net58);
INTERCONNECT SplitCLK_2_40_SplitCLK_6_35(net59_c1,net59);
INTERCONNECT SplitCLK_2_40_SplitCLK_4_39(net60_c1,net60);
INTERCONNECT SplitCLK_4_39_SplitCLK_2_37(net61_c1,net61);
INTERCONNECT SplitCLK_4_39_SplitCLK_6_38(net62_c1,net62);
INTERCONNECT SplitCLK_6_38_SplitCLK_2_42(net63_c1,net63);
INTERCONNECT SplitCLK_6_38_SplitCLK_4_50(net64_c1,net64);
INTERCONNECT SplitCLK_2_37_SplitCLK_2_51(net65_c1,net65);
INTERCONNECT SplitCLK_2_37_SplitCLK_4_36(net66_c1,net66);
INTERCONNECT SplitCLK_4_36_DFFT_24__FPB_n51(net67_c1,net67);
INTERCONNECT SplitCLK_4_36_DFFT_28__FPB_n55(net68_c1,net68);
INTERCONNECT SplitCLK_6_35_SplitCLK_4_33(net69_c1,net69);
INTERCONNECT SplitCLK_6_35_SplitCLK_6_34(net70_c1,net70);
INTERCONNECT SplitCLK_6_34_SplitCLK_2_43(net71_c1,net71);
INTERCONNECT SplitCLK_6_34_SplitCLK_4_47(net72_c1,net72);
INTERCONNECT SplitCLK_4_33_SplitCLK_2_49(net73_c1,net73);
INTERCONNECT SplitCLK_4_33_SplitCLK_4_32(net74_c1,net74);
INTERCONNECT SplitCLK_4_32_XOR2T_11_n11(net75_c1,net75);
INTERCONNECT SplitCLK_4_32_DFFT_26__FPB_n53(net76_c1,net76);
INTERCONNECT SplitCLK_0_31_SplitCLK_6_26(net77_c1,net77);
INTERCONNECT SplitCLK_0_31_SplitCLK_4_30(net78_c1,net78);
INTERCONNECT SplitCLK_4_30_SplitCLK_4_28(net79_c1,net79);
INTERCONNECT SplitCLK_4_30_SplitCLK_2_29(net80_c1,net80);
INTERCONNECT SplitCLK_2_29_SplitCLK_2_45(net81_c1,net81);
INTERCONNECT SplitCLK_2_29_SplitCLK_4_46(net82_c1,net82);
INTERCONNECT SplitCLK_4_28_SplitCLK_2_48(net83_c1,net83);
INTERCONNECT SplitCLK_4_28_SplitCLK_4_27(net84_c1,net84);
INTERCONNECT SplitCLK_4_27_XOR2T_10_n10(net85_c1,net85);
INTERCONNECT SplitCLK_4_27_XOR2T_15_sum1(net86_c1,net86);
INTERCONNECT SplitCLK_6_26_SplitCLK_4_23(net87_c1,net87);
INTERCONNECT SplitCLK_6_26_SplitCLK_2_25(net88_c1,net88);
INTERCONNECT SplitCLK_2_25_SplitCLK_4_41(net89_c1,net89);
INTERCONNECT SplitCLK_2_25_SplitCLK_4_24(net90_c1,net90);
INTERCONNECT SplitCLK_4_24_AND2T_13_n13(net91_c1,net91);
INTERCONNECT SplitCLK_4_24_AND2T_17_n17(net92_c1,net92);
INTERCONNECT SplitCLK_4_23_SplitCLK_4_44(net93_c1,net93);
INTERCONNECT SplitCLK_4_23_SplitCLK_4_22(net94_c1,net94);
INTERCONNECT SplitCLK_4_22_XOR2T_9_n9(net95_c1,net95);
INTERCONNECT SplitCLK_4_22_DFFT_22__FPB_n49(net96_c1,net96);
INTERCONNECT GCLK_Pad_SplitCLK_0_52(GCLK_Pad,net97);

endmodule
