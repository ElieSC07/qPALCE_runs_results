`timescale 1ps / 1fs
module tb;
	reg GCLK_Pad;
	reg a0_Pad;
	reg a1_Pad;
	reg b0_Pad;
	reg a2_Pad;
	reg b1_Pad;
	reg a3_Pad;
	reg b2_Pad;
	reg b3_Pad;
	reg cin_Pad;
	wire cout_Pad;
	wire sum0_Pad;
	wire sum1_Pad;
	wire sum2_Pad;
	wire sum3_Pad;
	KSA4_route topLevel(.GCLK_Pad(GCLK_Pad), .a0_Pad(a0_Pad), .a1_Pad(a1_Pad), .b0_Pad(b0_Pad), .a2_Pad(a2_Pad), .b1_Pad(b1_Pad), .a3_Pad(a3_Pad), .b2_Pad(b2_Pad), .b3_Pad(b3_Pad), .cin_Pad(cin_Pad), .cout_Pad(cout_Pad), .sum0_Pad(sum0_Pad), .sum1_Pad(sum1_Pad), .sum2_Pad(sum2_Pad), .sum3_Pad(sum3_Pad));
	initial begin
		$dumpfile("KSA4_route.vcd");
		$dumpvars(0,tb);
		$sdf_annotate("KSA4_route_qVsim.sdf");
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#40;
		a0_Pad = 1'd1;
		a1_Pad = 1'd1;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd1;
		a3_Pad = 1'd0;
		b2_Pad = 1'd1;
		b3_Pad = 1'd1;
		cin_Pad = 1'd1;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd1;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd0;
		a1_Pad = 1'd1;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd1;
		b2_Pad = 1'd1;
		b3_Pad = 1'd1;
		cin_Pad = 1'd1;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd1;
		a1_Pad = 1'd0;
		b0_Pad = 1'd1;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd1;
		b3_Pad = 1'd0;
		cin_Pad = 1'd1;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd1;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd1;
		b1_Pad = 1'd1;
		a3_Pad = 1'd0;
		b2_Pad = 1'd1;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd1;
		a2_Pad = 1'd0;
		b1_Pad = 1'd1;
		a3_Pad = 1'd1;
		b2_Pad = 1'd1;
		b3_Pad = 1'd1;
		cin_Pad = 1'd0;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd1;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd1;
		a1_Pad = 1'd1;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd1;
		a3_Pad = 1'd1;
		b2_Pad = 1'd1;
		b3_Pad = 1'd1;
		cin_Pad = 1'd0;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd1;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd1;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd0;
		a1_Pad = 1'd1;
		b0_Pad = 1'd0;
		a2_Pad = 1'd1;
		b1_Pad = 1'd0;
		a3_Pad = 1'd1;
		b2_Pad = 1'd1;
		b3_Pad = 1'd1;
		cin_Pad = 1'd1;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#38;
		a0_Pad = 1'd1;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd1;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd1;
		#2;
		a0_Pad = 1'd0;
		a1_Pad = 1'd0;
		b0_Pad = 1'd0;
		a2_Pad = 1'd0;
		b1_Pad = 1'd0;
		a3_Pad = 1'd0;
		b2_Pad = 1'd0;
		b3_Pad = 1'd0;
		cin_Pad = 1'd0;
		#38;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#78;
		GCLK_Pad = 1;
		#2;
		GCLK_Pad = 0;
		#10 $finish;
	end
endmodule
