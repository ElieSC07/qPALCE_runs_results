module TAP_route(
input GCLK_Pad,
input TMS_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output state_obs2_Pad,
output state_obs3_Pad);

wire TMS_Pad;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire TRST_Pad;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire state_obs0_Pad;
wire net405_c1;
wire state_obs1_Pad;
wire net406_c1;
wire state_obs2_Pad;
wire net407_c1;
wire state_obs3_Pad;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire net486_c1;
wire net486;
wire net487_c1;
wire net487;
wire net488_c1;
wire net488;
wire net489_c1;
wire net489;
wire net490_c1;
wire net490;
wire net491_c1;
wire net491;
wire net492_c1;
wire net492;
wire net493_c1;
wire net493;
wire net494_c1;
wire net494;
wire net495_c1;
wire net495;
wire net496_c1;
wire net496;
wire net497_c1;
wire net497;
wire net498_c1;
wire net498;
wire net499_c1;
wire net499;
wire net500_c1;
wire net500;
wire net501_c1;
wire net501;
wire net502_c1;
wire net502;
wire net503_c1;
wire net503;
wire net504_c1;
wire net504;
wire net505_c1;
wire net505;
wire net506_c1;
wire net506;
wire net507_c1;
wire net507;
wire net508_c1;
wire net508;
wire net509_c1;
wire net509;
wire net510_c1;
wire net510;
wire net511_c1;
wire net511;
wire net512_c1;
wire net512;
wire net513_c1;
wire net513;
wire net514_c1;
wire net514;
wire net515_c1;
wire net515;
wire net516_c1;
wire net516;
wire net517_c1;
wire net517;
wire net518_c1;
wire net518;
wire net519_c1;
wire net519;
wire net520_c1;
wire net520;
wire net521_c1;
wire net521;
wire net522_c1;
wire net522;
wire net523_c1;
wire net523;
wire net524_c1;
wire net524;
wire net525_c1;
wire net525;
wire net526_c1;
wire net526;
wire net527_c1;
wire net527;
wire net528_c1;
wire net528;
wire net529_c1;
wire net529;
wire net530_c1;
wire net530;
wire net531_c1;
wire net531;
wire net532_c1;
wire net532;
wire net533_c1;
wire net533;
wire net534_c1;
wire net534;
wire net535_c1;
wire net535;
wire net536_c1;
wire net536;
wire net537_c1;
wire net537;
wire net538_c1;
wire net538;
wire net539_c1;
wire net539;
wire net540_c1;
wire net540;
wire net541_c1;
wire net541;
wire net542_c1;
wire net542;
wire net543_c1;
wire net543;
wire net544_c1;
wire net544;
wire net545_c1;
wire net545;
wire net546_c1;
wire net546;
wire net547_c1;
wire net547;
wire net548_c1;
wire net548;
wire net549_c1;
wire net549;
wire net550_c1;
wire net550;
wire net551_c1;
wire net551;
wire net552_c1;
wire net552;
wire net553_c1;
wire net553;
wire net554_c1;
wire net554;
wire net555_c1;
wire net555;
wire net556_c1;
wire net556;
wire net557_c1;
wire net557;
wire net558_c1;
wire net558;
wire net559_c1;
wire net559;
wire net560_c1;
wire net560;
wire net561_c1;
wire net561;
wire net562_c1;
wire net562;
wire net563_c1;
wire net563;
wire net564_c1;
wire net564;
wire net565_c1;
wire net565;
wire net566_c1;
wire net566;
wire net567_c1;
wire net567;
wire net568_c1;
wire net568;
wire net569_c1;
wire net569;
wire net570_c1;
wire net570;
wire net571_c1;
wire net571;
wire net572_c1;
wire net572;
wire net573_c1;
wire net573;
wire net574_c1;
wire net574;
wire net575_c1;
wire net575;
wire net576_c1;
wire net576;
wire net577_c1;
wire net577;
wire net578_c1;
wire net578;
wire net579_c1;
wire net579;
wire net580_c1;
wire net580;
wire net581_c1;
wire net581;
wire net582_c1;
wire net582;
wire net583_c1;
wire net583;
wire net584_c1;
wire net584;
wire net585_c1;
wire net585;
wire net586_c1;
wire net586;
wire net587_c1;
wire net587;
wire net588_c1;
wire net588;
wire net589_c1;
wire net589;
wire net590_c1;
wire net590;
wire net591_c1;
wire net591;
wire net592_c1;
wire net592;
wire net593_c1;
wire net593;
wire net594_c1;
wire net594;
wire net595_c1;
wire net595;
wire net596_c1;
wire net596;
wire net597_c1;
wire net597;
wire net598_c1;
wire net598;
wire net599_c1;
wire net599;
wire net600_c1;
wire net600;
wire net601_c1;
wire net601;
wire net602_c1;
wire net602;
wire net603_c1;
wire net603;
wire net604_c1;
wire net604;
wire net605_c1;
wire net605;
wire net606_c1;
wire net606;
wire net607_c1;
wire net607;
wire net608_c1;
wire net608;
wire net609_c1;
wire net609;
wire net610_c1;
wire net610;
wire net611_c1;
wire net611;
wire net612_c1;
wire net612;
wire net613_c1;
wire net613;
wire net614_c1;
wire net614;
wire net615_c1;
wire net615;
wire net616_c1;
wire net616;
wire net617_c1;
wire net617;
wire net618_c1;
wire net618;
wire net619_c1;
wire net619;
wire net620_c1;
wire net620;
wire net621_c1;
wire net621;
wire net622_c1;
wire net622;
wire net623_c1;
wire net623;
wire net624_c1;
wire net624;
wire net625_c1;
wire net625;
wire net626_c1;
wire net626;
wire net627_c1;
wire net627;
wire net628_c1;
wire net628;
wire net629_c1;
wire net629;
wire net630_c1;
wire net630;
wire net631_c1;
wire net631;
wire net632_c1;
wire net632;
wire net633_c1;
wire net633;
wire net634_c1;
wire net634;
wire net635_c1;
wire net635;
wire net636_c1;
wire net636;
wire net637_c1;
wire net637;
wire net638_c1;
wire net638;
wire net639_c1;
wire net639;
wire net640_c1;
wire net640;
wire net641_c1;
wire net641;
wire net642_c1;
wire net642;
wire net643_c1;
wire net643;
wire net644_c1;
wire net644;
wire net645_c1;
wire net645;
wire net646_c1;
wire net646;
wire net647_c1;
wire net647;
wire net648_c1;
wire net648;
wire net649_c1;
wire net649;
wire net650_c1;
wire net650;
wire net651_c1;
wire net651;
wire net652_c1;
wire net652;
wire net653_c1;
wire net653;
wire net654_c1;
wire net654;
wire net655_c1;
wire net655;
wire net656_c1;
wire net656;
wire net657_c1;
wire net657;
wire net658_c1;
wire net658;
wire net659_c1;
wire net659;
wire net660_c1;
wire net660;
wire net661_c1;
wire net661;
wire net662_c1;
wire net662;
wire net663_c1;
wire net663;
wire net664_c1;
wire net664;
wire net665_c1;
wire net665;
wire net666_c1;
wire net666;
wire net667_c1;
wire net667;
wire net668_c1;
wire net668;
wire net669_c1;
wire net669;
wire net670_c1;
wire net670;
wire net671_c1;
wire net671;
wire net672_c1;
wire net672;
wire net673_c1;
wire net673;
wire net674_c1;
wire net674;
wire net675_c1;
wire net675;
wire net676_c1;
wire net676;
wire net677_c1;
wire net677;
wire net678_c1;
wire net678;
wire net679_c1;
wire net679;
wire net680_c1;
wire net680;
wire net681_c1;
wire net681;
wire net682_c1;
wire net682;
wire net683_c1;
wire net683;
wire net684_c1;
wire net684;
wire net685_c1;
wire net685;
wire net686_c1;
wire net686;
wire net687_c1;
wire net687;
wire net688_c1;
wire net688;
wire net689_c1;
wire net689;
wire net690_c1;
wire net690;
wire net691_c1;
wire net691;
wire net692_c1;
wire net692;
wire net693_c1;
wire net693;
wire net694_c1;
wire net694;
wire net695_c1;
wire net695;
wire net696_c1;
wire net696;
wire net697_c1;
wire net697;
wire net698_c1;
wire net698;
wire net699_c1;
wire net699;
wire net700_c1;
wire net700;
wire net701_c1;
wire net701;
wire net702_c1;
wire net702;
wire net703_c1;
wire net703;
wire net704_c1;
wire net704;
wire net705_c1;
wire net705;
wire net706_c1;
wire net706;
wire net707_c1;
wire net707;
wire net708_c1;
wire net708;
wire net709_c1;
wire net709;
wire net710_c1;
wire net710;
wire net711_c1;
wire net711;
wire net712_c1;
wire net712;
wire net713_c1;
wire net713;
wire net714_c1;
wire net714;
wire net715_c1;
wire net715;
wire net716_c1;
wire net716;
wire net717_c1;
wire net717;
wire net718_c1;
wire net718;
wire net719_c1;
wire net719;
wire net720_c1;
wire net720;
wire net721_c1;
wire net721;
wire net722_c1;
wire net722;
wire net723_c1;
wire net723;
wire net724_c1;
wire net724;
wire net725_c1;
wire net725;
wire net726_c1;
wire net726;
wire net727_c1;
wire net727;
wire net728_c1;
wire net728;
wire net729_c1;
wire net729;
wire net730_c1;
wire net730;
wire net731_c1;
wire net731;
wire net732_c1;
wire net732;
wire net733_c1;
wire net733;
wire net734_c1;
wire net734;
wire net735_c1;
wire net735;
wire net736_c1;
wire net736;
wire net737_c1;
wire net737;
wire net738_c1;
wire net738;
wire net739_c1;
wire net739;
wire net740_c1;
wire net740;
wire net741_c1;
wire net741;
wire net742_c1;
wire net742;
wire net743_c1;
wire net743;
wire net744_c1;
wire net744;
wire net745_c1;
wire net745;
wire net746_c1;
wire net746;
wire net747_c1;
wire net747;
wire net748_c1;
wire net748;
wire net749_c1;
wire net749;
wire net750_c1;
wire net750;
wire net751_c1;
wire net751;
wire net752_c1;
wire net752;
wire net753_c1;
wire net753;
wire net754_c1;
wire net754;
wire net755_c1;
wire net755;
wire net756_c1;
wire net756;
wire net757_c1;
wire net757;
wire net758_c1;
wire net758;
wire net759_c1;
wire net759;
wire net760_c1;
wire net760;
wire net761_c1;
wire net761;
wire net762_c1;
wire net762;
wire net763_c1;
wire net763;
wire net764_c1;
wire net764;
wire net765_c1;
wire net765;
wire net766_c1;
wire net766;
wire net767_c1;
wire net767;
wire net768_c1;
wire net768;
wire net769_c1;
wire net769;
wire net770_c1;
wire net770;
wire net771_c1;
wire net771;
wire net772_c1;
wire net772;
wire net773_c1;
wire net773;
wire net774_c1;
wire net774;
wire net775_c1;
wire net775;
wire net776_c1;
wire net776;
wire net777_c1;
wire net777;
wire net778_c1;
wire net778;
wire net779_c1;
wire net779;
wire net780_c1;
wire net780;
wire net781_c1;
wire net781;
wire net782_c1;
wire net782;
wire net783_c1;
wire net783;
wire net784_c1;
wire net784;
wire net785_c1;
wire net785;
wire net786_c1;
wire net786;
wire net787_c1;
wire net787;
wire net788_c1;
wire net788;
wire net789_c1;
wire net789;
wire net790_c1;
wire net790;
wire net791_c1;
wire net791;
wire net792_c1;
wire net792;
wire net793_c1;
wire net793;
wire net794_c1;
wire net794;
wire net795_c1;
wire net795;
wire net796_c1;
wire net796;
wire net797_c1;
wire net797;
wire net798_c1;
wire net798;
wire net799_c1;
wire net799;
wire net800_c1;
wire net800;
wire net801_c1;
wire net801;
wire net802_c1;
wire net802;
wire net803_c1;
wire net803;
wire net804_c1;
wire net804;
wire net805_c1;
wire net805;
wire net806_c1;
wire net806;
wire net807_c1;
wire net807;
wire net808_c1;
wire net808;
wire net809_c1;
wire net809;
wire net810_c1;
wire net810;
wire net811_c1;
wire net811;
wire net812_c1;
wire net812;
wire net813_c1;
wire net813;
wire net814_c1;
wire net814;
wire net815_c1;
wire net815;
wire net816_c1;
wire net816;
wire net817_c1;
wire net817;
wire net818_c1;
wire net818;
wire net819_c1;
wire net819;
wire net820_c1;
wire net820;
wire net821_c1;
wire net821;
wire net822_c1;
wire net822;
wire net823_c1;
wire net823;
wire net824_c1;
wire net824;
wire net825_c1;
wire net825;
wire net826_c1;
wire net826;
wire net827_c1;
wire net827;
wire net828_c1;
wire net828;
wire net829_c1;
wire net829;
wire net830_c1;
wire net830;
wire net831_c1;
wire net831;
wire net832_c1;
wire net832;
wire net833_c1;
wire net833;
wire net834_c1;
wire net834;
wire net835_c1;
wire net835;
wire net836_c1;
wire net836;
wire net837_c1;
wire net837;
wire net838_c1;
wire net838;
wire net839_c1;
wire net839;
wire net840_c1;
wire net840;
wire net841_c1;
wire net841;
wire net842_c1;
wire net842;
wire net843_c1;
wire net843;
wire net844_c1;
wire net844;
wire net845_c1;
wire net845;
wire net846_c1;
wire net846;
wire net847_c1;
wire net847;
wire net848_c1;
wire net848;
wire net849_c1;
wire net849;
wire net850_c1;
wire net850;
wire net851_c1;
wire net851;
wire net852_c1;
wire net852;
wire net853_c1;
wire net853;
wire net854_c1;
wire net854;
wire net855_c1;
wire net855;
wire net856_c1;
wire net856;
wire net857_c1;
wire net857;
wire net858_c1;
wire net858;
wire net859_c1;
wire net859;
wire net860_c1;
wire net860;
wire net861_c1;
wire net861;
wire net862_c1;
wire net862;
wire net863_c1;
wire net863;
wire net864_c1;
wire net864;
wire net865_c1;
wire net865;
wire net866_c1;
wire net866;
wire net867_c1;
wire net867;
wire net868_c1;
wire net868;
wire net869_c1;
wire net869;
wire net870_c1;
wire net870;
wire net871_c1;
wire net871;
wire net872_c1;
wire net872;
wire net873_c1;
wire net873;
wire net874_c1;
wire net874;
wire net875_c1;
wire net875;
wire net876_c1;
wire net876;
wire net877_c1;
wire net877;
wire net878_c1;
wire net878;
wire net879_c1;
wire net879;
wire net880_c1;
wire net880;
wire net881_c1;
wire net881;
wire net882_c1;
wire net882;
wire net883_c1;
wire net883;
wire net884_c1;
wire net884;
wire net885_c1;
wire net885;
wire net886_c1;
wire net886;
wire net887_c1;
wire net887;
wire net888_c1;
wire net888;
wire net889_c1;
wire net889;
wire net890_c1;
wire net890;
wire net891_c1;
wire net891;
wire net892_c1;
wire net892;
wire net893_c1;
wire net893;
wire net894_c1;
wire net894;
wire net895_c1;
wire net895;
wire net896_c1;
wire net896;
wire net897_c1;
wire net897;
wire net898_c1;
wire net898;
wire net899_c1;
wire net899;
wire net900_c1;
wire net900;
wire net901_c1;
wire net901;
wire GCLK_Pad;
wire net902;
wire net903_c1;
wire net903;
wire net904_c1;
wire net904;
wire net905_c1;
wire net905;
wire net906_c1;
wire net906;
wire net907_c1;
wire net907;
wire net908_c1;
wire net908;
wire net909_c1;
wire net909;
wire net910_c1;
wire net910;

DFFT DFFT_199__FPB_n619(net748,net327,net336_c1);
DFFT DFFT_245_state_obs3(net826,net378,net407_c1);
AND2T AND2T_103_n139(net782,net279,net148,net94_c1);
DFFT DFFT_239_state_obs2(net662,net391,net406_c1);
NOTT NOTT_8_n32(net429,net111,net2_c1);
NOTT NOTT_9_n33(net480,net200,net4_c1);
AND2T AND2T_20_n44(net812,net136,net120,net13_c1);
AND2T AND2T_12_n36(net572,net195,net217,net14_c1);
AND2T AND2T_21_n45(net894,net167,net152,net17_c1);
AND2T AND2T_22_n46(net724,net224,net255,net22_c1);
AND2T AND2T_14_n38(net814,net208,net349,net23_c1);
AND2T AND2T_31_n55(net630,net228,net233,net26_c1);
AND2T AND2T_15_n39(net616,net250,net227,net28_c1);
AND2T AND2T_40_n64(net636,net25,net168,net31_c1);
AND2T AND2T_32_n56(net806,net163,net323,net32_c1);
AND2T AND2T_17_n41(net856,net223,net125,net3_c1);
AND2T AND2T_25_n49(net428,net258,net341,net38_c1);
AND2T AND2T_26_n50(net427,net151,net348,net5_c1);
AND2T AND2T_18_n42(net558,net110,net359,net6_c1);
AND2T AND2T_42_n66(net822,net257,net384,net42_c1);
AND2T AND2T_34_n58(net488,net48,net21,net43_c1);
AND2T AND2T_27_n51(net870,net141,net358,net8_c1);
AND2T AND2T_19_n43(net794,net246,net234,net9_c1);
AND2T AND2T_43_n67(net578,net264,net166,net47_c1);
AND2T AND2T_36_n60(net576,net135,net357,net11_c1);
AND2T AND2T_28_n52(net631,net262,net146,net12_c1);
AND2T AND2T_44_n68(net489,net181,net332,net52_c1);
AND2T AND2T_37_n61(net634,net216,net226,net15_c1);
AND2T AND2T_61_n85(net468,net4,net383,net54_c1);
AND2T AND2T_53_n77(net469,net51,net345,net55_c1);
AND2T AND2T_45_n69(net617,net150,net339,net56_c1);
AND2T AND2T_46_n70(net798,net213,net189,net19_c1);
AND2T AND2T_38_n62(net620,net252,net910,net20_c1);
AND2T AND2T_70_n94(net482,net53,net289,net57_c1);
AND2T AND2T_62_n86(net823,net254,net390,net58_c1);
AND2T AND2T_47_n71(net637,net19,net179,net24_c1);
AND2T AND2T_39_n63(net799,net202,net377,net25_c1);
AND2T AND2T_71_n95(net768,net114,net292,net60_c1);
AND2T AND2T_63_n87(net880,net58,net197,net61_c1);
AND2T AND2T_56_n80(net526,net62,net394,net29_c1);
AND2T AND2T_72_n96(net852,net103,net214,net63_c1);
AND2T AND2T_64_n88(net644,net199,net393,net64_c1);
AND2T AND2T_57_n81(net628,net178,net240,net34_c1);
AND2T AND2T_65_n89(net656,net64,net263,net66_c1);
AND2T AND2T_59_n83(net426,net190,net401,net45_c1);
AND2T AND2T_75_n99(net516,net69,net287,net68_c1);
OR2T OR2T_30_n54(net708,net241,net315,net21_c1);
OR2T OR2T_23_n47(net546,net9,net301,net27_c1);
OR2T OR2T_24_n48(net544,net27,net307,net33_c1);
OR2T OR2T_41_n65(net622,net31,net20,net36_c1);
OR2T OR2T_33_n57(net486,net247,net340,net37_c1);
OR2T OR2T_50_n74(net474,net35,net346,net41_c1);
OR2T OR2T_51_n75(net475,net41,net43,net46_c1);
OR2T OR2T_35_n59(net472,net37,net347,net48_c1);
OR2T OR2T_60_n84(net623,net261,net367,net50_c1);
OR2T OR2T_52_n76(net532,net46,net356,net51_c1);
OR2T OR2T_29_n53(net808,net12,net5,net16_c1);
OR2T OR2T_54_n78(net533,net96,net162,net59_c1);
OR2T OR2T_55_n79(net538,net174,net355,net62_c1);
OR2T OR2T_48_n72(net425,net183,net182,net30_c1);
OR2T OR2T_49_n73(net573,net30,net52,net35_c1);
OR2T OR2T_73_n97(net858,net63,net295,net65_c1);
OR2T OR2T_66_n90(net635,net201,net397,net39_c1);
OR2T OR2T_58_n82(net795,net34,net98,net40_c1);
OR2T OR2T_74_n98(net780,net60,net300,net67_c1);
OR2T OR2T_67_n91(net629,net39,net50,net44_c1);
OR2T OR2T_68_n92(net539,net44,net399,net49_c1);
OR2T OR2T_69_n93(net527,net49,net29,net53_c1);
DFFT DFFT_106__PIPL_n154(net600,net408,net266_c1);
DFFT DFFT_107__PIPL_n155(net664,net409,net267_c1);
DFFT DFFT_108__PIPL_n156(net828,net90,net268_c1);
NOTT NOTT_10_n34(net857,net205,net7_c1);
NOTT NOTT_11_n35(net813,net221,net10_c1);
NOTT NOTT_13_n37(net884,net237,net18_c1);
NOTT NOTT_16_n40(net842,net253,net1_c1);
DFFT DFFT_109__PIPL_n157(net892,net75,net269_c1);
DFFT DFFT_97_state0_buf(net598,net225,net408_c1);
AND2T AND2T_83_n107(net746,net81,net293,net83_c1);
AND2T AND2T_84_n108(net762,net106,net314,net85_c1);
AND2T AND2T_77_n101(net684,net68,net67,net70_c1);
AND2T AND2T_85_n109(net725,net171,net220,net87_c1);
AND2T AND2T_86_n110(net774,net87,net235,net71_c1);
AND2T AND2T_78_n102(net809,net130,net129,net72_c1);
AND2T AND2T_94_n118(net694,net86,net338,net88_c1);
AND2T AND2T_87_n111(net872,net905,net906,net73_c1);
AND2T AND2T_79_n103(net807,net72,net299,net74_c1);
AND2T AND2T_89_n113(net834,net259,net239,net78_c1);
DFFT DFFT_110__FBL_n530(net424,net187,net270_c1);
DFFT DFFT_111__FBL_n531(net658,net184,net271_c1);
DFFT DFFT_120__FBL_n540(net895,net330,net272_c1);
DFFT DFFT_112__FBL_n532(net696,net298,net273_c1);
DFFT DFFT_104__FPB_n152(net458,net155,net282_c1);
DFFT DFFT_200__FPB_n620(net754,net336,net290_c1);
DFFT DFFT_121__FBL_n541(net423,net337,net274_c1);
DFFT DFFT_113__FBL_n533(net460,net305,net275_c1);
DFFT DFFT_98_state1_buf(net827,net230,net409_c1);
DFFT DFFT_105__FPB_n153(net446,net232,net283_c1);
DFFT DFFT_201__FPB_n621(net749,net290,net293_c1);
DFFT DFFT_114__FBL_n534(net562,net102,net276_c1);
DFFT DFFT_210__FPB_n630(net690,net128,net296_c1);
DFFT DFFT_202__FPB_n622(net776,net134,net297_c1);
DFFT DFFT_130__FPB_n550(net709,net22,net301_c1);
DFFT DFFT_122__FPB_n542(net738,net188,net298_c1);
DFFT DFFT_115__FBL_n535(net601,net97,net277_c1);
DFFT DFFT_211__FPB_n631(net422,net296,net302_c1);
DFFT DFFT_203__FPB_n623(net775,net297,net303_c1);
DFFT DFFT_131__FPB_n551(net421,net28,net307_c1);
DFFT DFFT_123__FPB_n543(net454,net194,net305_c1);
DFFT DFFT_116__FBL_n536(net752,net313,net278_c1);
DFFT DFFT_220__FPB_n640(net586,net372,net308_c1);
DFFT DFFT_212__FPB_n632(net678,net302,net309_c1);
DFFT DFFT_204__FPB_n624(net763,net303,net314_c1);
DFFT DFFT_140__FPB_n560(net710,net376,net315_c1);
DFFT DFFT_132__FPB_n552(net704,net119,net312_c1);
DFFT DFFT_124__FPB_n544(net740,net101,net313_c1);
DFFT DFFT_117__FBL_n537(net777,net321,net279_c1);
DFFT DFFT_221__FPB_n641(net592,net308,net316_c1);
DFFT DFFT_213__FPB_n633(net679,net309,net317_c1);
DFFT DFFT_205__FPB_n625(net866,net143,net322_c1);
DFFT DFFT_141__FPB_n561(net722,net140,net323_c1);
DFFT DFFT_133__FPB_n553(net705,net312,net320_c1);
DFFT DFFT_125__FPB_n545(net755,net108,net321_c1);
DFFT DFFT_118__FBL_n538(net564,net185,net280_c1);
DFFT DFFT_230__FPB_n650(net648,net386,net324_c1);
DFFT DFFT_222__FPB_n642(net604,net907,net325_c1);
DFFT DFFT_214__FPB_n634(net691,net317,net326_c1);
DFFT DFFT_206__FPB_n626(net836,net78,net331_c1);
DFFT DFFT_150__FPB_n570(net530,net389,net332_c1);
DFFT DFFT_142__FPB_n562(net487,net115,net328_c1);
DFFT DFFT_134__FPB_n554(net540,net320,net329_c1);
DFFT DFFT_126__FPB_n546(net753,net186,net330_c1);
DFFT DFFT_119__FBL_n539(net565,net206,net281_c1);
DFFT DFFT_231__FPB_n651(net650,net324,net333_c1);
DFFT DFFT_223__FPB_n643(net590,net325,net334_c1);
DFFT DFFT_215__FPB_n635(net697,net326,net338_c1);
DFFT DFFT_207__FPB_n627(net769,net71,net335_c1);
DFFT DFFT_151__FPB_n571(net864,net229,net339_c1);
DFFT DFFT_143__FPB_n563(net531,net328,net340_c1);
DFFT DFFT_135__FPB_n555(net541,net329,net341_c1);
DFFT DFFT_127__FPB_n547(net741,net191,net337_c1);
OR2T OR2T_80_n104(net800,net74,net95,net77_c1);
OR2T OR2T_81_n105(net711,net77,net158,net79_c1);
OR2T OR2T_90_n114(net873,net73,net331,net80_c1);
OR2T OR2T_82_n106(net695,net70,net306,net81_c1);
OR2T OR2T_91_n115(net871,net80,net118,net82_c1);
OR2T OR2T_76_n100(net510,net193,net294,net69_c1);
OR2T OR2T_92_n116(net766,net82,net344,net84_c1);
OR2T OR2T_93_n117(net718,net84,net354,net86_c1);
DFFT DFFT_240__FPB_n660(net886,net269,net342_c1);
DFFT DFFT_216__FPB_n636(net893,net909,net343_c1);
DFFT DFFT_208__FPB_n628(net767,net335,net344_c1);
DFFT DFFT_160__FPB_n580(net448,net396,net345_c1);
DFFT DFFT_152__FPB_n572(net570,net176,net346_c1);
DFFT DFFT_144__FPB_n564(net571,net26,net347_c1);
DFFT DFFT_136__FPB_n556(net853,net251,net348_c1);
DFFT DFFT_128__FPB_n548(net659,net131,net349_c1);
OR2T OR2T_96_n120(net887,net170,net343,net75_c1);
OR2T OR2T_88_n112(net865,net218,net7,net76_c1);
DFFT DFFT_241__FPB_n661(net898,net342,net350_c1);
DFFT DFFT_233__FPB_n653(net829,net268,net351_c1);
DFFT DFFT_225__FPB_n645(net657,net267,net352_c1);
DFFT DFFT_217__FPB_n637(net606,net266,net353_c1);
DFFT DFFT_209__FPB_n629(net739,net85,net354_c1);
DFFT DFFT_161__FPB_n581(net545,net59,net355_c1);
DFFT DFFT_153__FPB_n573(net547,net38,net356_c1);
DFFT DFFT_145__FPB_n565(net837,net154,net357_c1);
DFFT DFFT_137__FPB_n557(net881,net243,net358_c1);
DFFT DFFT_129__FPB_n549(net559,net210,net359_c1);
DFFT DFFT_242__FPB_n662(net899,net350,net360_c1);
DFFT DFFT_234__FPB_n654(net840,net351,net361_c1);
DFFT DFFT_226__FPB_n646(net420,net352,net362_c1);
DFFT DFFT_218__FPB_n638(net593,net353,net363_c1);
DFFT DFFT_170__FPB_n590(net621,net265,net367_c1);
DFFT DFFT_162__FPB_n582(net419,net117,net364_c1);
DFFT DFFT_154__FPB_n574(net512,net249,net365_c1);
DFFT DFFT_146__FPB_n566(net579,net172,net368_c1);
DFFT DFFT_138__FPB_n558(net716,net207,net366_c1);
DFFT DFFT_243__FPB_n663(net900,net360,net369_c1);
DFFT DFFT_235__FPB_n655(net843,net361,net370_c1);
DFFT DFFT_227__FPB_n647(net649,net362,net371_c1);
DFFT DFFT_219__FPB_n639(net587,net363,net372_c1);
DFFT DFFT_171__FPB_n591(net418,net123,net373_c1);
DFFT DFFT_163__FPB_n583(net461,net364,net374_c1);
DFFT DFFT_155__FPB_n575(net417,net365,net375_c1);
DFFT DFFT_147__FPB_n567(net801,net139,net377_c1);
DFFT DFFT_139__FPB_n559(net717,net366,net376_c1);
DFFT DFFT_180__FPB_n600(net498,net403,net284_c1);
DFFT DFFT_244__FPB_n664(net901,net369,net378_c1);
DFFT DFFT_236__FPB_n656(net885,net370,net379_c1);
DFFT DFFT_228__FPB_n648(net651,net371,net380_c1);
DFFT DFFT_172__FPB_n592(net473,net373,net383_c1);
DFFT DFFT_164__FPB_n584(net416,net374,net381_c1);
DFFT DFFT_156__FPB_n576(net442,net375,net382_c1);
DFFT DFFT_148__FPB_n568(net415,net144,net384_c1);
DFFT DFFT_181__FPB_n601(net414,net284,net285_c1);
DFFT DFFT_237__FPB_n657(net663,net379,net385_c1);
DFFT DFFT_229__FPB_n649(net607,net380,net386_c1);
DFFT DFFT_173__FPB_n593(net835,net113,net390_c1);
DFFT DFFT_165__FPB_n585(net504,net381,net387_c1);
DFFT DFFT_157__FPB_n577(net443,net382,net388_c1);
DFFT DFFT_149__FPB_n569(net481,net204,net389_c1);
DFFT DFFT_190__FPB_n610(net518,net319,net287_c1);
DFFT DFFT_182__FPB_n602(net455,net285,net286_c1);
DFFT DFFT_238__FPB_n658(net665,net385,net391_c1);
DFFT DFFT_174__FPB_n594(net577,net138,net393_c1);
DFFT DFFT_166__FPB_n586(net483,net387,net394_c1);
DFFT DFFT_158__FPB_n578(net413,net388,net392_c1);
SPLITT Split_300_n720(net127,net103_c1,net189_c1);
SPLITT Split_301_n721(net92,net104_c1,net192_c1);
SPLITT Split_302_n722(net192,net110_c1,net195_c1);
SPLITT Split_310_n730(net282,net107_c1,net196_c1);
SPLITT Split_303_n723(net104,net113_c1,net199_c1);
SPLITT Split_311_n731(net196,net115_c1,net200_c1);
SPLITT Split_304_n724(net93,net116_c1,net203_c1);
SPLITT Split_312_n732(net107,net117_c1,net204_c1);
SPLITT Split_320_n740(net242,net120_c1,net205_c1);
SPLITT Split_305_n725(net203,net125_c1,net208_c1);
SPLITT Split_313_n733(net283,net121_c1,net209_c1);
SPLITT Split_321_n741(net153,net123_c1,net210_c1);
SPLITT Split_250_n670(net161,net128_c1,net212_c1);
SPLITT Split_306_n726(net116,net130_c1,net213_c1);
SPLITT Split_314_n734(net209,net129_c1,net214_c1);
SPLITT Split_322_n742(net281,net126_c1,net215_c1);
SPLITT Split_330_n750(net159,net131_c1,net216_c1);
SPLITT Split_251_n671(net10,net133_c1,net218_c1);
SPLITT Split_307_n727(net94,net132_c1,net219_c1);
SPLITT Split_315_n735(net121,net134_c1,net220_c1);
SPLITT Split_323_n743(net215,net136_c1,net221_c1);
SPLITT Split_252_n672(net14,net137_c1,net222_c1);
SPLITT Split_260_n680(net173,net141_c1,net223_c1);
SPLITT Split_308_n728(net219,net140_c1,net224_c1);
SPLITT Split_316_n736(net270,net138_c1,net225_c1);
SPLITT Split_324_n744(net126,net139_c1,net226_c1);
SPLITT Split_253_n673(net222,net146_c1,net227_c1);
SPLITT Split_261_n681(net3,net145_c1,net228_c1);
SPLITT Split_309_n729(net132,net143_c1,net229_c1);
SPLITT Split_317_n737(net271,net144_c1,net230_c1);
SPLITT Split_325_n745(net272,net142_c1,net231_c1);
SPLITT Split_246_n666(net0,net147_c1,net232_c1);
SPLITT Split_254_n674(net137,net150_c1,net233_c1);
SPLITT Split_262_n682(net145,net151_c1,net234_c1);
SPLITT Split_270_n690(net175,net149_c1,net235_c1);
SPLITT Split_318_n738(net278,net148_c1,net236_c1);
SPLITT Split_326_n746(net231,net152_c1,net237_c1);
SPLITT Split_247_n667(net147,net155_c1,net238_c1);
SPLITT Split_255_n675(net18,net156_c1,net239_c1);
SPLITT Split_263_n683(net6,net157_c1,net240_c1);
SPLITT Split_271_n691(net16,net158_c1,net241_c1);
SPLITT Split_319_n739(net280,net153_c1,net242_c1);
SPLITT Split_327_n747(net142,net154_c1,net243_c1);
SPLITT Split_280_n700(net180,net95_c1,net181_c1);
SPLITT Split_248_n668(net2,net161_c1,net244_c1);
SPLITT Split_256_n676(net23,net160_c1,net245_c1);
SPLITT Split_264_n684(net157,net163_c1,net246_c1);
SPLITT Split_272_n692(net32,net162_c1,net247_c1);
SPLITT Split_328_n748(net274,net159_c1,net248_c1);
SPLITT Split_281_n701(net56,net96_c1,net182_c1);
SPLITT Split_249_n669(net244,net164_c1,net249_c1);
SPLITT Split_257_n677(net245,net168_c1,net250_c1);
SPLITT Split_265_n685(net13,net165_c1,net251_c1);
SPLITT Split_273_n693(net11,net166_c1,net252_c1);
SPLITT Split_329_n749(net248,net167_c1,net253_c1);
DFFT DFFT_191__FPB_n611(net502,net275,net288_c1);
DFFT DFFT_183__FPB_n603(net449,net286,net289_c1);
SPLITT Split_282_n702(net24,net98_c1,net183_c1);
SPLITT Split_290_n710(net124,net97_c1,net184_c1);
DFFT DFFT_175__FPB_n595(net645,net66,net397_c1);
DFFT DFFT_167__FPB_n587(net517,net122,net395_c1);
DFFT DFFT_159__FPB_n579(net447,net392,net396_c1);
SPLITT Split_258_n678(net160,net170_c1,net254_c1);
SPLITT Split_266_n686(net165,net171_c1,net255_c1);
SPLITT Split_274_n694(net15,net169_c1,net256_c1);
SPLITT Split_283_n703(net55,net100_c1,net185_c1);
SPLITT Split_291_n711(net83,net99_c1,net186_c1);
SPLITT Split_259_n679(net1,net173_c1,net257_c1);
SPLITT Split_267_n687(net33,net174_c1,net258_c1);
SPLITT Split_275_n695(net169,net172_c1,net259_c1);
SPLITT Split_284_n704(net100,net102_c1,net187_c1);
SPLITT Split_292_n712(net99,net101_c1,net188_c1);
SPLITT Split_268_n688(net8,net175_c1,net260_c1);
SPLITT Split_276_n696(net36,net176_c1,net261_c1);
SPLITT Split_285_n705(net40,net106_c1,net190_c1);
SPLITT Split_293_n713(net88,net105_c1,net191_c1);
SPLITT Split_269_n689(net260,net178_c1,net262_c1);
SPLITT Split_277_n697(net42,net177_c1,net263_c1);
SPLITT Split_286_n706(net54,net109_c1,net193_c1);
SPLITT Split_294_n714(net105,net108_c1,net194_c1);
SPLITT Split_278_n698(net177,net179_c1,net264_c1);
SPLITT Split_287_n707(net109,net114_c1,net197_c1);
SPLITT Split_295_n715(net89,net112_c1,net198_c1);
SPLITT Split_279_n699(net47,net180_c1,net265_c1);
SPLITT Split_288_n708(net61,net118_c1,net201_c1);
SPLITT Split_296_n716(net198,net119_c1,net202_c1);
SPLITT Split_289_n709(net57,net124_c1,net206_c1);
SPLITT Split_297_n717(net112,net122_c1,net207_c1);
SPLITT Split_298_n718(net91,net127_c1,net211_c1);
SPLITT Split_299_n719(net211,net135_c1,net217_c1);
NOTT NOTT_100_n136(net563,net276,net91_c1);
NOTT NOTT_101_n137(net599,net908,net92_c1);
NOTT NOTT_102_n138(net867,net236,net93_c1);
DFFT DFFT_192__FPB_n612(net503,net288,net291_c1);
DFFT DFFT_184__FPB_n604(net783,net149,net292_c1);
DFFT DFFT_176__FPB_n596(net719,net45,net399_c1);
DFFT DFFT_168__FPB_n588(net519,net395,net398_c1);
DFFT DFFT_193__FPB_n613(net505,net291,net294_c1);
DFFT DFFT_185__FPB_n605(net859,net133,net295_c1);
DFFT DFFT_177__FPB_n597(net513,net164,net400_c1);
DFFT DFFT_169__FPB_n589(net682,net904,net401_c1);
DFFT DFFT_194__FPB_n614(net815,net256,net299_c1);
DFFT DFFT_186__FPB_n606(net781,net65,net300_c1);
DFFT DFFT_178__FPB_n598(net511,net400,net402_c1);
DFFT DFFT_195__FPB_n615(net723,net79,net306_c1);
DFFT DFFT_187__FPB_n607(net685,net273,net304_c1);
DFFT DFFT_179__FPB_n599(net499,net402,net403_c1);
DFFT DFFT_196__FPB_n616(net734,net212,net310_c1);
DFFT DFFT_188__FPB_n608(net683,net903,net311_c1);
NOTT NOTT_95_n119(net841,net156,net90_c1);
NOTT NOTT_99_n135(net459,net238,net89_c1);
DFFT DFFT_197__FPB_n617(net735,net310,net318_c1);
DFFT DFFT_189__FPB_n609(net412,net311,net319_c1);
DFFT DFFT_224_state_obs0(net591,net334,net404_c1);
DFFT DFFT_232_state_obs1(net605,net333,net405_c1);
DFFT DFFT_198__FPB_n618(net747,net318,net327_c1);
SPLITT SplitCLK_4_239(net896,net900_c1,net901_c1);
SPLITT SplitCLK_4_240(net897,net898_c1,net899_c1);
SPLITT SplitCLK_6_241(net888,net896_c1,net897_c1);
SPLITT SplitCLK_4_242(net890,net895_c1,net894_c1);
SPLITT SplitCLK_0_243(net891,net892_c1,net893_c1);
SPLITT SplitCLK_2_244(net889,net890_c1,net891_c1);
SPLITT SplitCLK_4_245(net874,net889_c1,net888_c1);
SPLITT SplitCLK_4_246(net882,net886_c1,net887_c1);
SPLITT SplitCLK_4_247(net883,net884_c1,net885_c1);
SPLITT SplitCLK_6_248(net876,net882_c1,net883_c1);
SPLITT SplitCLK_4_249(net879,net881_c1,net880_c1);
SPLITT SplitCLK_2_250(net877,net878_c1,net879_c1);
SPLITT SplitCLK_2_251(net875,net877_c1,net876_c1);
SPLITT SplitCLK_6_252(net844,net874_c1,net875_c1);
SPLITT SplitCLK_4_253(net868,net872_c1,net873_c1);
SPLITT SplitCLK_4_254(net869,net870_c1,net871_c1);
SPLITT SplitCLK_6_255(net860,net868_c1,net869_c1);
SPLITT SplitCLK_4_256(net862,net866_c1,net867_c1);
SPLITT SplitCLK_4_257(net863,net865_c1,net864_c1);
SPLITT SplitCLK_4_258(net861,net863_c1,net862_c1);
SPLITT SplitCLK_0_259(net846,net860_c1,net861_c1);
SPLITT SplitCLK_4_260(net854,net858_c1,net859_c1);
SPLITT SplitCLK_4_261(net855,net856_c1,net857_c1);
SPLITT SplitCLK_6_262(net848,net854_c1,net855_c1);
SPLITT SplitCLK_4_263(net851,net852_c1,net853_c1);
SPLITT SplitCLK_2_264(net849,net850_c1,net851_c1);
SPLITT SplitCLK_2_265(net847,net849_c1,net848_c1);
SPLITT SplitCLK_4_266(net845,net847_c1,net846_c1);
SPLITT SplitCLK_0_267(net784,net844_c1,net845_c1);
SPLITT SplitCLK_4_268(net838,net842_c1,net843_c1);
SPLITT SplitCLK_4_269(net839,net841_c1,net840_c1);
SPLITT SplitCLK_6_270(net830,net838_c1,net839_c1);
SPLITT SplitCLK_4_271(net832,net836_c1,net837_c1);
SPLITT SplitCLK_4_272(net833,net834_c1,net835_c1);
SPLITT SplitCLK_4_273(net831,net833_c1,net832_c1);
SPLITT SplitCLK_4_274(net816,net831_c1,net830_c1);
SPLITT SplitCLK_4_275(net824,net829_c1,net828_c1);
SPLITT SplitCLK_4_276(net825,net826_c1,net827_c1);
SPLITT SplitCLK_6_277(net818,net824_c1,net825_c1);
SPLITT SplitCLK_4_278(net821,net823_c1,net822_c1);
SPLITT SplitCLK_2_279(net819,net820_c1,net821_c1);
SPLITT SplitCLK_6_280(net817,net819_c1,net818_c1);
SPLITT SplitCLK_6_281(net786,net816_c1,net817_c1);
SPLITT SplitCLK_0_282(net810,net814_c1,net815_c1);
SPLITT SplitCLK_4_283(net811,net812_c1,net813_c1);
SPLITT SplitCLK_4_284(net802,net811_c1,net810_c1);
SPLITT SplitCLK_4_285(net804,net809_c1,net808_c1);
SPLITT SplitCLK_4_286(net805,net807_c1,net806_c1);
SPLITT SplitCLK_4_287(net803,net805_c1,net804_c1);
SPLITT SplitCLK_0_288(net788,net802_c1,net803_c1);
SPLITT SplitCLK_4_289(net796,net800_c1,net801_c1);
SPLITT SplitCLK_4_290(net797,net798_c1,net799_c1);
SPLITT SplitCLK_6_291(net790,net796_c1,net797_c1);
SPLITT SplitCLK_4_292(net793,net795_c1,net794_c1);
SPLITT SplitCLK_4_293(net791,net792_c1,net793_c1);
SPLITT SplitCLK_4_294(net789,net791_c1,net790_c1);
SPLITT SplitCLK_4_295(net787,net789_c1,net788_c1);
SPLITT SplitCLK_2_296(net785,net787_c1,net786_c1);
SPLITT SplitCLK_6_297(net666,net784_c1,net785_c1);
SPLITT SplitCLK_4_298(net778,net783_c1,net782_c1);
SPLITT SplitCLK_0_299(net779,net781_c1,net780_c1);
SPLITT SplitCLK_0_300(net770,net779_c1,net778_c1);
SPLITT SplitCLK_4_301(net772,net776_c1,net777_c1);
SPLITT SplitCLK_4_302(net773,net775_c1,net774_c1);
SPLITT SplitCLK_4_303(net771,net773_c1,net772_c1);
SPLITT SplitCLK_4_304(net756,net770_c1,net771_c1);
SPLITT SplitCLK_4_305(net764,net768_c1,net769_c1);
SPLITT SplitCLK_4_306(net765,net766_c1,net767_c1);
SPLITT SplitCLK_6_307(net758,net764_c1,net765_c1);
SPLITT SplitCLK_4_308(net761,net762_c1,net763_c1);
SPLITT SplitCLK_6_309(net759,net761_c1,net760_c1);
SPLITT SplitCLK_4_310(net757,net759_c1,net758_c1);
SPLITT SplitCLK_6_311(net726,net756_c1,net757_c1);
SPLITT SplitCLK_4_312(net750,net755_c1,net754_c1);
SPLITT SplitCLK_0_313(net751,net752_c1,net753_c1);
SPLITT SplitCLK_0_314(net742,net751_c1,net750_c1);
SPLITT SplitCLK_4_315(net744,net748_c1,net749_c1);
SPLITT SplitCLK_4_316(net745,net747_c1,net746_c1);
SPLITT SplitCLK_6_317(net743,net744_c1,net745_c1);
SPLITT SplitCLK_4_318(net728,net743_c1,net742_c1);
SPLITT SplitCLK_4_319(net736,net741_c1,net740_c1);
SPLITT SplitCLK_0_320(net737,net739_c1,net738_c1);
SPLITT SplitCLK_6_321(net730,net736_c1,net737_c1);
SPLITT SplitCLK_4_322(net733,net734_c1,net735_c1);
SPLITT SplitCLK_4_323(net731,net732_c1,net733_c1);
SPLITT SplitCLK_2_324(net729,net731_c1,net730_c1);
SPLITT SplitCLK_4_325(net727,net729_c1,net728_c1);
SPLITT SplitCLK_0_326(net668,net726_c1,net727_c1);
SPLITT SplitCLK_4_327(net720,net725_c1,net724_c1);
SPLITT SplitCLK_4_328(net721,net723_c1,net722_c1);
SPLITT SplitCLK_4_329(net712,net721_c1,net720_c1);
SPLITT SplitCLK_4_330(net714,net718_c1,net719_c1);
SPLITT SplitCLK_4_331(net715,net717_c1,net716_c1);
SPLITT SplitCLK_4_332(net713,net715_c1,net714_c1);
SPLITT SplitCLK_0_333(net698,net712_c1,net713_c1);
SPLITT SplitCLK_4_334(net706,net710_c1,net711_c1);
SPLITT SplitCLK_4_335(net707,net709_c1,net708_c1);
SPLITT SplitCLK_6_336(net700,net706_c1,net707_c1);
SPLITT SplitCLK_4_337(net703,net705_c1,net704_c1);
SPLITT SplitCLK_2_338(net701,net703_c1,net702_c1);
SPLITT SplitCLK_6_339(net699,net700_c1,net701_c1);
SPLITT SplitCLK_6_340(net670,net698_c1,net699_c1);
SPLITT SplitCLK_4_341(net692,net697_c1,net696_c1);
SPLITT SplitCLK_0_342(net693,net694_c1,net695_c1);
SPLITT SplitCLK_0_343(net686,net693_c1,net692_c1);
SPLITT SplitCLK_4_344(net689,net691_c1,net690_c1);
SPLITT SplitCLK_2_345(net687,net688_c1,net689_c1);
SPLITT SplitCLK_4_346(net672,net687_c1,net686_c1);
SPLITT SplitCLK_4_347(net680,net684_c1,net685_c1);
SPLITT SplitCLK_0_348(net681,net682_c1,net683_c1);
SPLITT SplitCLK_6_349(net674,net680_c1,net681_c1);
SPLITT SplitCLK_4_350(net677,net679_c1,net678_c1);
SPLITT SplitCLK_4_351(net675,net676_c1,net677_c1);
SPLITT SplitCLK_2_352(net673,net674_c1,net675_c1);
SPLITT SplitCLK_4_353(net671,net673_c1,net672_c1);
SPLITT SplitCLK_2_354(net669,net671_c1,net670_c1);
SPLITT SplitCLK_4_355(net667,net669_c1,net668_c1);
SPLITT SplitCLK_0_356(net410,net666_c1,net667_c1);
SPLITT SplitCLK_4_357(net660,net664_c1,net665_c1);
SPLITT SplitCLK_0_358(net661,net662_c1,net663_c1);
SPLITT SplitCLK_6_359(net652,net660_c1,net661_c1);
SPLITT SplitCLK_4_360(net654,net659_c1,net658_c1);
SPLITT SplitCLK_4_361(net655,net656_c1,net657_c1);
SPLITT SplitCLK_4_362(net653,net655_c1,net654_c1);
SPLITT SplitCLK_0_363(net638,net652_c1,net653_c1);
SPLITT SplitCLK_4_364(net646,net650_c1,net651_c1);
SPLITT SplitCLK_4_365(net647,net648_c1,net649_c1);
SPLITT SplitCLK_6_366(net640,net646_c1,net647_c1);
SPLITT SplitCLK_4_367(net643,net645_c1,net644_c1);
SPLITT SplitCLK_6_368(net641,net643_c1,net642_c1);
SPLITT SplitCLK_6_369(net639,net640_c1,net641_c1);
SPLITT SplitCLK_6_370(net608,net638_c1,net639_c1);
SPLITT SplitCLK_4_371(net632,net637_c1,net636_c1);
SPLITT SplitCLK_4_372(net633,net634_c1,net635_c1);
SPLITT SplitCLK_6_373(net624,net632_c1,net633_c1);
SPLITT SplitCLK_4_374(net626,net630_c1,net631_c1);
SPLITT SplitCLK_4_375(net627,net629_c1,net628_c1);
SPLITT SplitCLK_4_376(net625,net627_c1,net626_c1);
SPLITT SplitCLK_0_377(net610,net624_c1,net625_c1);
SPLITT SplitCLK_4_378(net618,net623_c1,net622_c1);
SPLITT SplitCLK_0_379(net619,net620_c1,net621_c1);
SPLITT SplitCLK_6_380(net612,net618_c1,net619_c1);
SPLITT SplitCLK_4_381(net615,net616_c1,net617_c1);
SPLITT SplitCLK_4_382(net613,net614_c1,net615_c1);
SPLITT SplitCLK_4_383(net611,net612_c1,net613_c1);
SPLITT SplitCLK_4_384(net609,net611_c1,net610_c1);
SPLITT SplitCLK_6_385(net548,net608_c1,net609_c1);
SPLITT SplitCLK_4_386(net602,net606_c1,net607_c1);
SPLITT SplitCLK_0_387(net603,net604_c1,net605_c1);
SPLITT SplitCLK_0_388(net594,net603_c1,net602_c1);
SPLITT SplitCLK_4_389(net596,net600_c1,net601_c1);
SPLITT SplitCLK_4_390(net597,net598_c1,net599_c1);
SPLITT SplitCLK_4_391(net595,net597_c1,net596_c1);
SPLITT SplitCLK_4_392(net580,net594_c1,net595_c1);
SPLITT SplitCLK_4_393(net588,net592_c1,net593_c1);
SPLITT SplitCLK_0_394(net589,net590_c1,net591_c1);
SPLITT SplitCLK_0_395(net582,net589_c1,net588_c1);
SPLITT SplitCLK_4_396(net585,net587_c1,net586_c1);
SPLITT SplitCLK_6_397(net583,net585_c1,net584_c1);
SPLITT SplitCLK_2_398(net581,net582_c1,net583_c1);
SPLITT SplitCLK_6_399(net550,net580_c1,net581_c1);
SPLITT SplitCLK_4_400(net574,net579_c1,net578_c1);
SPLITT SplitCLK_0_401(net575,net577_c1,net576_c1);
SPLITT SplitCLK_6_402(net566,net574_c1,net575_c1);
SPLITT SplitCLK_4_403(net568,net572_c1,net573_c1);
SPLITT SplitCLK_4_404(net569,net571_c1,net570_c1);
SPLITT SplitCLK_4_405(net567,net569_c1,net568_c1);
SPLITT SplitCLK_0_406(net552,net566_c1,net567_c1);
SPLITT SplitCLK_4_407(net560,net564_c1,net565_c1);
SPLITT SplitCLK_4_408(net561,net562_c1,net563_c1);
SPLITT SplitCLK_2_409(net554,net560_c1,net561_c1);
SPLITT SplitCLK_4_410(net557,net559_c1,net558_c1);
SPLITT SplitCLK_4_411(net555,net556_c1,net557_c1);
SPLITT SplitCLK_2_412(net553,net555_c1,net554_c1);
SPLITT SplitCLK_4_413(net551,net553_c1,net552_c1);
SPLITT SplitCLK_2_414(net549,net551_c1,net550_c1);
SPLITT SplitCLK_6_415(net430,net548_c1,net549_c1);
SPLITT SplitCLK_4_416(net542,net547_c1,net546_c1);
SPLITT SplitCLK_4_417(net543,net545_c1,net544_c1);
SPLITT SplitCLK_6_418(net534,net542_c1,net543_c1);
SPLITT SplitCLK_4_419(net536,net541_c1,net540_c1);
SPLITT SplitCLK_4_420(net537,net539_c1,net538_c1);
SPLITT SplitCLK_4_421(net535,net537_c1,net536_c1);
SPLITT SplitCLK_6_422(net520,net535_c1,net534_c1);
SPLITT SplitCLK_4_423(net528,net533_c1,net532_c1);
SPLITT SplitCLK_4_424(net529,net531_c1,net530_c1);
SPLITT SplitCLK_6_425(net522,net528_c1,net529_c1);
SPLITT SplitCLK_4_426(net525,net526_c1,net527_c1);
SPLITT SplitCLK_6_427(net523,net525_c1,net524_c1);
SPLITT SplitCLK_6_428(net521,net522_c1,net523_c1);
SPLITT SplitCLK_4_429(net490,net521_c1,net520_c1);
SPLITT SplitCLK_4_430(net514,net519_c1,net518_c1);
SPLITT SplitCLK_4_431(net515,net517_c1,net516_c1);
SPLITT SplitCLK_4_432(net506,net515_c1,net514_c1);
SPLITT SplitCLK_4_433(net508,net513_c1,net512_c1);
SPLITT SplitCLK_2_434(net509,net511_c1,net510_c1);
SPLITT SplitCLK_4_435(net507,net509_c1,net508_c1);
SPLITT SplitCLK_0_436(net492,net506_c1,net507_c1);
SPLITT SplitCLK_4_437(net500,net504_c1,net505_c1);
SPLITT SplitCLK_4_438(net501,net502_c1,net503_c1);
SPLITT SplitCLK_4_439(net494,net501_c1,net500_c1);
SPLITT SplitCLK_4_440(net497,net498_c1,net499_c1);
SPLITT SplitCLK_4_441(net495,net496_c1,net497_c1);
SPLITT SplitCLK_6_442(net493,net494_c1,net495_c1);
SPLITT SplitCLK_4_443(net491,net493_c1,net492_c1);
SPLITT SplitCLK_0_444(net432,net490_c1,net491_c1);
SPLITT SplitCLK_4_445(net484,net489_c1,net488_c1);
SPLITT SplitCLK_4_446(net485,net486_c1,net487_c1);
SPLITT SplitCLK_6_447(net476,net484_c1,net485_c1);
SPLITT SplitCLK_4_448(net478,net482_c1,net483_c1);
SPLITT SplitCLK_4_449(net479,net481_c1,net480_c1);
SPLITT SplitCLK_2_450(net477,net478_c1,net479_c1);
SPLITT SplitCLK_4_451(net462,net477_c1,net476_c1);
SPLITT SplitCLK_4_452(net470,net474_c1,net475_c1);
SPLITT SplitCLK_4_453(net471,net473_c1,net472_c1);
SPLITT SplitCLK_2_454(net464,net470_c1,net471_c1);
SPLITT SplitCLK_4_455(net467,net469_c1,net468_c1);
SPLITT SplitCLK_6_456(net465,net467_c1,net466_c1);
SPLITT SplitCLK_6_457(net463,net464_c1,net465_c1);
SPLITT SplitCLK_6_458(net434,net462_c1,net463_c1);
SPLITT SplitCLK_4_459(net456,net460_c1,net461_c1);
SPLITT SplitCLK_4_460(net457,net458_c1,net459_c1);
SPLITT SplitCLK_6_461(net450,net456_c1,net457_c1);
SPLITT SplitCLK_4_462(net453,net454_c1,net455_c1);
SPLITT SplitCLK_2_463(net451,net452_c1,net453_c1);
SPLITT SplitCLK_0_464(net436,net450_c1,net451_c1);
SPLITT SplitCLK_4_465(net444,net448_c1,net449_c1);
SPLITT SplitCLK_4_466(net445,net447_c1,net446_c1);
SPLITT SplitCLK_6_467(net438,net444_c1,net445_c1);
SPLITT SplitCLK_4_468(net441,net443_c1,net442_c1);
SPLITT SplitCLK_4_469(net439,net440_c1,net441_c1);
SPLITT SplitCLK_2_470(net437,net439_c1,net438_c1);
SPLITT SplitCLK_4_471(net435,net437_c1,net436_c1);
SPLITT SplitCLK_2_472(net433,net435_c1,net434_c1);
SPLITT SplitCLK_4_473(net431,net433_c1,net432_c1);
SPLITT SplitCLK_2_474(net411,net431_c1,net430_c1);
wire dummy0;
SPLITT SplitCLK_2_475(net732,net429_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_2_476(net702,net428_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_477(net850,net427_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_478(net760,net426_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_479(net614,net425_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_4_480(net584,net424_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_2_481(net878,net423_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_2_482(net688,net422_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_2_483(net792,net421_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_2_484(net642,net420_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_4_485(net466,net419_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_4_486(net556,net418_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_2_487(net452,net417_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_4_488(net524,net416_c1,dummy13);
wire dummy14;
SPLITT SplitCLK_2_489(net820,net415_c1,dummy14);
wire dummy15;
SPLITT SplitCLK_2_490(net496,net414_c1,dummy15);
wire dummy16;
SPLITT SplitCLK_2_491(net440,net413_c1,dummy16);
wire dummy17;
SPLITT SplitCLK_2_492(net676,net412_c1,dummy17);
SPLITT SplitCLK_0_493(net902,net410_c1,net411_c1);
wire dummy18;
SPLITT Split_HOLD_586(net304,dummy18,net903_c1);
wire dummy19;
SPLITT Split_HOLD_587(net398,dummy19,net904_c1);
wire dummy20;
SPLITT Split_HOLD_588(net76,dummy20,net905_c1);
wire dummy21;
SPLITT Split_HOLD_589(net322,dummy21,net906_c1);
wire dummy22;
SPLITT Split_HOLD_590(net316,dummy22,net907_c1);
wire dummy23;
SPLITT Split_HOLD_591(net277,dummy23,net908_c1);
wire dummy24;
SPLITT Split_HOLD_592(net17,dummy24,net909_c1);
wire dummy25;
SPLITT Split_HOLD_593(net368,dummy25,net910_c1);
INTERCONNECT TMS_Pad_Split_246_n666(TMS_Pad,net0);
INTERCONNECT NOTT_16_n40_Split_259_n679(net1_c1,net1);
INTERCONNECT NOTT_8_n32_Split_248_n668(net2_c1,net2);
INTERCONNECT AND2T_17_n41_Split_261_n681(net3_c1,net3);
INTERCONNECT NOTT_9_n33_AND2T_61_n85(net4_c1,net4);
INTERCONNECT AND2T_26_n50_OR2T_29_n53(net5_c1,net5);
INTERCONNECT AND2T_18_n42_Split_263_n683(net6_c1,net6);
INTERCONNECT NOTT_10_n34_OR2T_88_n112(net7_c1,net7);
INTERCONNECT AND2T_27_n51_Split_268_n688(net8_c1,net8);
INTERCONNECT AND2T_19_n43_OR2T_23_n47(net9_c1,net9);
INTERCONNECT NOTT_11_n35_Split_251_n671(net10_c1,net10);
INTERCONNECT AND2T_36_n60_Split_273_n693(net11_c1,net11);
INTERCONNECT AND2T_28_n52_OR2T_29_n53(net12_c1,net12);
INTERCONNECT AND2T_20_n44_Split_265_n685(net13_c1,net13);
INTERCONNECT AND2T_12_n36_Split_252_n672(net14_c1,net14);
INTERCONNECT AND2T_37_n61_Split_274_n694(net15_c1,net15);
INTERCONNECT OR2T_29_n53_Split_271_n691(net16_c1,net16);
INTERCONNECT AND2T_21_n45_Split_HOLD_592(net17_c1,net17);
INTERCONNECT NOTT_13_n37_Split_255_n675(net18_c1,net18);
INTERCONNECT AND2T_46_n70_AND2T_47_n71(net19_c1,net19);
INTERCONNECT AND2T_38_n62_OR2T_41_n65(net20_c1,net20);
INTERCONNECT OR2T_30_n54_AND2T_34_n58(net21_c1,net21);
INTERCONNECT AND2T_22_n46_DFFT_130__FPB_n550(net22_c1,net22);
INTERCONNECT AND2T_14_n38_Split_256_n676(net23_c1,net23);
INTERCONNECT AND2T_47_n71_Split_282_n702(net24_c1,net24);
INTERCONNECT AND2T_39_n63_AND2T_40_n64(net25_c1,net25);
INTERCONNECT AND2T_31_n55_DFFT_144__FPB_n564(net26_c1,net26);
INTERCONNECT OR2T_23_n47_OR2T_24_n48(net27_c1,net27);
INTERCONNECT AND2T_15_n39_DFFT_131__FPB_n551(net28_c1,net28);
INTERCONNECT AND2T_56_n80_OR2T_69_n93(net29_c1,net29);
INTERCONNECT OR2T_48_n72_OR2T_49_n73(net30_c1,net30);
INTERCONNECT AND2T_40_n64_OR2T_41_n65(net31_c1,net31);
INTERCONNECT AND2T_32_n56_Split_272_n692(net32_c1,net32);
INTERCONNECT OR2T_24_n48_Split_267_n687(net33_c1,net33);
INTERCONNECT AND2T_57_n81_OR2T_58_n82(net34_c1,net34);
INTERCONNECT OR2T_49_n73_OR2T_50_n74(net35_c1,net35);
INTERCONNECT OR2T_41_n65_Split_276_n696(net36_c1,net36);
INTERCONNECT OR2T_33_n57_OR2T_35_n59(net37_c1,net37);
INTERCONNECT AND2T_25_n49_DFFT_153__FPB_n573(net38_c1,net38);
INTERCONNECT OR2T_66_n90_OR2T_67_n91(net39_c1,net39);
INTERCONNECT OR2T_58_n82_Split_285_n705(net40_c1,net40);
INTERCONNECT OR2T_50_n74_OR2T_51_n75(net41_c1,net41);
INTERCONNECT AND2T_42_n66_Split_277_n697(net42_c1,net42);
INTERCONNECT AND2T_34_n58_OR2T_51_n75(net43_c1,net43);
INTERCONNECT OR2T_67_n91_OR2T_68_n92(net44_c1,net44);
INTERCONNECT AND2T_59_n83_DFFT_176__FPB_n596(net45_c1,net45);
INTERCONNECT OR2T_51_n75_OR2T_52_n76(net46_c1,net46);
INTERCONNECT AND2T_43_n67_Split_279_n699(net47_c1,net47);
INTERCONNECT OR2T_35_n59_AND2T_34_n58(net48_c1,net48);
INTERCONNECT OR2T_68_n92_OR2T_69_n93(net49_c1,net49);
INTERCONNECT OR2T_60_n84_OR2T_67_n91(net50_c1,net50);
INTERCONNECT OR2T_52_n76_AND2T_53_n77(net51_c1,net51);
INTERCONNECT AND2T_44_n68_OR2T_49_n73(net52_c1,net52);
INTERCONNECT OR2T_69_n93_AND2T_70_n94(net53_c1,net53);
INTERCONNECT AND2T_61_n85_Split_286_n706(net54_c1,net54);
INTERCONNECT AND2T_53_n77_Split_283_n703(net55_c1,net55);
INTERCONNECT AND2T_45_n69_Split_281_n701(net56_c1,net56);
INTERCONNECT AND2T_70_n94_Split_289_n709(net57_c1,net57);
INTERCONNECT AND2T_62_n86_AND2T_63_n87(net58_c1,net58);
INTERCONNECT OR2T_54_n78_DFFT_161__FPB_n581(net59_c1,net59);
INTERCONNECT AND2T_71_n95_OR2T_74_n98(net60_c1,net60);
INTERCONNECT AND2T_63_n87_Split_288_n708(net61_c1,net61);
INTERCONNECT OR2T_55_n79_AND2T_56_n80(net62_c1,net62);
INTERCONNECT AND2T_72_n96_OR2T_73_n97(net63_c1,net63);
INTERCONNECT AND2T_64_n88_AND2T_65_n89(net64_c1,net64);
INTERCONNECT OR2T_73_n97_DFFT_186__FPB_n606(net65_c1,net65);
INTERCONNECT AND2T_65_n89_DFFT_175__FPB_n595(net66_c1,net66);
INTERCONNECT OR2T_74_n98_AND2T_77_n101(net67_c1,net67);
INTERCONNECT AND2T_75_n99_AND2T_77_n101(net68_c1,net68);
INTERCONNECT OR2T_76_n100_AND2T_75_n99(net69_c1,net69);
INTERCONNECT AND2T_77_n101_OR2T_82_n106(net70_c1,net70);
INTERCONNECT AND2T_86_n110_DFFT_207__FPB_n627(net71_c1,net71);
INTERCONNECT AND2T_78_n102_AND2T_79_n103(net72_c1,net72);
INTERCONNECT AND2T_87_n111_OR2T_90_n114(net73_c1,net73);
INTERCONNECT AND2T_79_n103_OR2T_80_n104(net74_c1,net74);
INTERCONNECT OR2T_96_n120_DFFT_109__PIPL_n157(net75_c1,net75);
INTERCONNECT OR2T_88_n112_Split_HOLD_588(net76_c1,net76);
INTERCONNECT OR2T_80_n104_OR2T_81_n105(net77_c1,net77);
INTERCONNECT AND2T_89_n113_DFFT_206__FPB_n626(net78_c1,net78);
INTERCONNECT OR2T_81_n105_DFFT_195__FPB_n615(net79_c1,net79);
INTERCONNECT OR2T_90_n114_OR2T_91_n115(net80_c1,net80);
INTERCONNECT OR2T_82_n106_AND2T_83_n107(net81_c1,net81);
INTERCONNECT OR2T_91_n115_OR2T_92_n116(net82_c1,net82);
INTERCONNECT AND2T_83_n107_Split_291_n711(net83_c1,net83);
INTERCONNECT OR2T_92_n116_OR2T_93_n117(net84_c1,net84);
INTERCONNECT AND2T_84_n108_DFFT_209__FPB_n629(net85_c1,net85);
INTERCONNECT OR2T_93_n117_AND2T_94_n118(net86_c1,net86);
INTERCONNECT AND2T_85_n109_AND2T_86_n110(net87_c1,net87);
INTERCONNECT AND2T_94_n118_Split_293_n713(net88_c1,net88);
INTERCONNECT NOTT_99_n135_Split_295_n715(net89_c1,net89);
INTERCONNECT NOTT_95_n119_DFFT_108__PIPL_n156(net90_c1,net90);
INTERCONNECT NOTT_100_n136_Split_298_n718(net91_c1,net91);
INTERCONNECT NOTT_101_n137_Split_301_n721(net92_c1,net92);
INTERCONNECT NOTT_102_n138_Split_304_n724(net93_c1,net93);
INTERCONNECT AND2T_103_n139_Split_307_n727(net94_c1,net94);
INTERCONNECT Split_280_n700_OR2T_80_n104(net95_c1,net95);
INTERCONNECT Split_281_n701_OR2T_54_n78(net96_c1,net96);
INTERCONNECT Split_290_n710_DFFT_115__FBL_n535(net97_c1,net97);
INTERCONNECT Split_282_n702_OR2T_58_n82(net98_c1,net98);
INTERCONNECT Split_291_n711_Split_292_n712(net99_c1,net99);
INTERCONNECT Split_283_n703_Split_284_n704(net100_c1,net100);
INTERCONNECT Split_292_n712_DFFT_124__FPB_n544(net101_c1,net101);
INTERCONNECT Split_284_n704_DFFT_114__FBL_n534(net102_c1,net102);
INTERCONNECT Split_300_n720_AND2T_72_n96(net103_c1,net103);
INTERCONNECT Split_301_n721_Split_303_n723(net104_c1,net104);
INTERCONNECT Split_293_n713_Split_294_n714(net105_c1,net105);
INTERCONNECT Split_285_n705_AND2T_84_n108(net106_c1,net106);
INTERCONNECT Split_310_n730_Split_312_n732(net107_c1,net107);
INTERCONNECT Split_294_n714_DFFT_125__FPB_n545(net108_c1,net108);
INTERCONNECT Split_286_n706_Split_287_n707(net109_c1,net109);
INTERCONNECT Split_302_n722_AND2T_18_n42(net110_c1,net110);
INTERCONNECT TRST_Pad_NOTT_8_n32(TRST_Pad,net111);
INTERCONNECT Split_295_n715_Split_297_n717(net112_c1,net112);
INTERCONNECT Split_303_n723_DFFT_173__FPB_n593(net113_c1,net113);
INTERCONNECT Split_287_n707_AND2T_71_n95(net114_c1,net114);
INTERCONNECT Split_311_n731_DFFT_142__FPB_n562(net115_c1,net115);
INTERCONNECT Split_304_n724_Split_306_n726(net116_c1,net116);
INTERCONNECT Split_312_n732_DFFT_162__FPB_n582(net117_c1,net117);
INTERCONNECT Split_288_n708_OR2T_91_n115(net118_c1,net118);
INTERCONNECT Split_296_n716_DFFT_132__FPB_n552(net119_c1,net119);
INTERCONNECT Split_320_n740_AND2T_20_n44(net120_c1,net120);
INTERCONNECT Split_313_n733_Split_315_n735(net121_c1,net121);
INTERCONNECT Split_297_n717_DFFT_167__FPB_n587(net122_c1,net122);
INTERCONNECT Split_321_n741_DFFT_171__FPB_n591(net123_c1,net123);
INTERCONNECT Split_289_n709_Split_290_n710(net124_c1,net124);
INTERCONNECT Split_305_n725_AND2T_17_n41(net125_c1,net125);
INTERCONNECT Split_322_n742_Split_324_n744(net126_c1,net126);
INTERCONNECT Split_298_n718_Split_300_n720(net127_c1,net127);
INTERCONNECT Split_250_n670_DFFT_210__FPB_n630(net128_c1,net128);
INTERCONNECT Split_314_n734_AND2T_78_n102(net129_c1,net129);
INTERCONNECT Split_306_n726_AND2T_78_n102(net130_c1,net130);
INTERCONNECT Split_330_n750_DFFT_128__FPB_n548(net131_c1,net131);
INTERCONNECT Split_307_n727_Split_309_n729(net132_c1,net132);
INTERCONNECT Split_251_n671_DFFT_185__FPB_n605(net133_c1,net133);
INTERCONNECT Split_315_n735_DFFT_202__FPB_n622(net134_c1,net134);
INTERCONNECT Split_299_n719_AND2T_36_n60(net135_c1,net135);
INTERCONNECT Split_323_n743_AND2T_20_n44(net136_c1,net136);
INTERCONNECT Split_252_n672_Split_254_n674(net137_c1,net137);
INTERCONNECT Split_316_n736_DFFT_174__FPB_n594(net138_c1,net138);
INTERCONNECT Split_324_n744_DFFT_147__FPB_n567(net139_c1,net139);
INTERCONNECT Split_308_n728_DFFT_141__FPB_n561(net140_c1,net140);
INTERCONNECT Split_260_n680_AND2T_27_n51(net141_c1,net141);
INTERCONNECT Split_325_n745_Split_327_n747(net142_c1,net142);
INTERCONNECT Split_309_n729_DFFT_205__FPB_n625(net143_c1,net143);
INTERCONNECT Split_317_n737_DFFT_148__FPB_n568(net144_c1,net144);
INTERCONNECT Split_261_n681_Split_262_n682(net145_c1,net145);
INTERCONNECT Split_253_n673_AND2T_28_n52(net146_c1,net146);
INTERCONNECT Split_246_n666_Split_247_n667(net147_c1,net147);
INTERCONNECT Split_318_n738_AND2T_103_n139(net148_c1,net148);
INTERCONNECT Split_270_n690_DFFT_184__FPB_n604(net149_c1,net149);
INTERCONNECT Split_254_n674_AND2T_45_n69(net150_c1,net150);
INTERCONNECT Split_262_n682_AND2T_26_n50(net151_c1,net151);
INTERCONNECT Split_326_n746_AND2T_21_n45(net152_c1,net152);
INTERCONNECT Split_319_n739_Split_321_n741(net153_c1,net153);
INTERCONNECT Split_327_n747_DFFT_145__FPB_n565(net154_c1,net154);
INTERCONNECT Split_247_n667_DFFT_104__FPB_n152(net155_c1,net155);
INTERCONNECT Split_255_n675_NOTT_95_n119(net156_c1,net156);
INTERCONNECT Split_263_n683_Split_264_n684(net157_c1,net157);
INTERCONNECT Split_271_n691_OR2T_81_n105(net158_c1,net158);
INTERCONNECT Split_328_n748_Split_330_n750(net159_c1,net159);
INTERCONNECT Split_256_n676_Split_258_n678(net160_c1,net160);
INTERCONNECT Split_248_n668_Split_250_n670(net161_c1,net161);
INTERCONNECT Split_272_n692_OR2T_54_n78(net162_c1,net162);
INTERCONNECT Split_264_n684_AND2T_32_n56(net163_c1,net163);
INTERCONNECT Split_249_n669_DFFT_177__FPB_n597(net164_c1,net164);
INTERCONNECT Split_265_n685_Split_266_n686(net165_c1,net165);
INTERCONNECT Split_273_n693_AND2T_43_n67(net166_c1,net166);
INTERCONNECT Split_329_n749_AND2T_21_n45(net167_c1,net167);
INTERCONNECT Split_257_n677_AND2T_40_n64(net168_c1,net168);
INTERCONNECT Split_274_n694_Split_275_n695(net169_c1,net169);
INTERCONNECT Split_258_n678_OR2T_96_n120(net170_c1,net170);
INTERCONNECT Split_266_n686_AND2T_85_n109(net171_c1,net171);
INTERCONNECT Split_275_n695_DFFT_146__FPB_n566(net172_c1,net172);
INTERCONNECT Split_259_n679_Split_260_n680(net173_c1,net173);
INTERCONNECT Split_267_n687_OR2T_55_n79(net174_c1,net174);
INTERCONNECT Split_268_n688_Split_270_n690(net175_c1,net175);
INTERCONNECT Split_276_n696_DFFT_152__FPB_n572(net176_c1,net176);
INTERCONNECT Split_277_n697_Split_278_n698(net177_c1,net177);
INTERCONNECT Split_269_n689_AND2T_57_n81(net178_c1,net178);
INTERCONNECT Split_278_n698_AND2T_47_n71(net179_c1,net179);
INTERCONNECT Split_279_n699_Split_280_n700(net180_c1,net180);
INTERCONNECT Split_280_n700_AND2T_44_n68(net181_c1,net181);
INTERCONNECT Split_281_n701_OR2T_48_n72(net182_c1,net182);
INTERCONNECT Split_282_n702_OR2T_48_n72(net183_c1,net183);
INTERCONNECT Split_290_n710_DFFT_111__FBL_n531(net184_c1,net184);
INTERCONNECT Split_283_n703_DFFT_118__FBL_n538(net185_c1,net185);
INTERCONNECT Split_291_n711_DFFT_126__FPB_n546(net186_c1,net186);
INTERCONNECT Split_284_n704_DFFT_110__FBL_n530(net187_c1,net187);
INTERCONNECT Split_292_n712_DFFT_122__FPB_n542(net188_c1,net188);
INTERCONNECT Split_300_n720_AND2T_46_n70(net189_c1,net189);
INTERCONNECT Split_285_n705_AND2T_59_n83(net190_c1,net190);
INTERCONNECT Split_293_n713_DFFT_127__FPB_n547(net191_c1,net191);
INTERCONNECT Split_301_n721_Split_302_n722(net192_c1,net192);
INTERCONNECT Split_286_n706_OR2T_76_n100(net193_c1,net193);
INTERCONNECT Split_294_n714_DFFT_123__FPB_n543(net194_c1,net194);
INTERCONNECT Split_302_n722_AND2T_12_n36(net195_c1,net195);
INTERCONNECT Split_310_n730_Split_311_n731(net196_c1,net196);
INTERCONNECT Split_287_n707_AND2T_63_n87(net197_c1,net197);
INTERCONNECT Split_295_n715_Split_296_n716(net198_c1,net198);
INTERCONNECT Split_303_n723_AND2T_64_n88(net199_c1,net199);
INTERCONNECT Split_311_n731_NOTT_9_n33(net200_c1,net200);
INTERCONNECT Split_288_n708_OR2T_66_n90(net201_c1,net201);
INTERCONNECT Split_296_n716_AND2T_39_n63(net202_c1,net202);
INTERCONNECT Split_304_n724_Split_305_n725(net203_c1,net203);
INTERCONNECT Split_312_n732_DFFT_149__FPB_n569(net204_c1,net204);
INTERCONNECT Split_320_n740_NOTT_10_n34(net205_c1,net205);
INTERCONNECT Split_289_n709_DFFT_119__FBL_n539(net206_c1,net206);
INTERCONNECT Split_297_n717_DFFT_138__FPB_n558(net207_c1,net207);
INTERCONNECT Split_305_n725_AND2T_14_n38(net208_c1,net208);
INTERCONNECT Split_313_n733_Split_314_n734(net209_c1,net209);
INTERCONNECT Split_321_n741_DFFT_129__FPB_n549(net210_c1,net210);
INTERCONNECT Split_298_n718_Split_299_n719(net211_c1,net211);
INTERCONNECT Split_250_n670_DFFT_196__FPB_n616(net212_c1,net212);
INTERCONNECT Split_306_n726_AND2T_46_n70(net213_c1,net213);
INTERCONNECT Split_314_n734_AND2T_72_n96(net214_c1,net214);
INTERCONNECT Split_322_n742_Split_323_n743(net215_c1,net215);
INTERCONNECT Split_330_n750_AND2T_37_n61(net216_c1,net216);
INTERCONNECT Split_299_n719_AND2T_12_n36(net217_c1,net217);
INTERCONNECT Split_251_n671_OR2T_88_n112(net218_c1,net218);
INTERCONNECT Split_307_n727_Split_308_n728(net219_c1,net219);
INTERCONNECT Split_315_n735_AND2T_85_n109(net220_c1,net220);
INTERCONNECT Split_323_n743_NOTT_11_n35(net221_c1,net221);
INTERCONNECT Split_252_n672_Split_253_n673(net222_c1,net222);
INTERCONNECT Split_260_n680_AND2T_17_n41(net223_c1,net223);
INTERCONNECT Split_308_n728_AND2T_22_n46(net224_c1,net224);
INTERCONNECT Split_316_n736_DFFT_97_state0_buf(net225_c1,net225);
INTERCONNECT Split_324_n744_AND2T_37_n61(net226_c1,net226);
INTERCONNECT Split_253_n673_AND2T_15_n39(net227_c1,net227);
INTERCONNECT Split_261_n681_AND2T_31_n55(net228_c1,net228);
INTERCONNECT Split_309_n729_DFFT_151__FPB_n571(net229_c1,net229);
INTERCONNECT Split_317_n737_DFFT_98_state1_buf(net230_c1,net230);
INTERCONNECT Split_325_n745_Split_326_n746(net231_c1,net231);
INTERCONNECT Split_246_n666_DFFT_105__FPB_n153(net232_c1,net232);
INTERCONNECT Split_254_n674_AND2T_31_n55(net233_c1,net233);
INTERCONNECT Split_262_n682_AND2T_19_n43(net234_c1,net234);
INTERCONNECT Split_270_n690_AND2T_86_n110(net235_c1,net235);
INTERCONNECT Split_318_n738_NOTT_102_n138(net236_c1,net236);
INTERCONNECT Split_326_n746_NOTT_13_n37(net237_c1,net237);
INTERCONNECT Split_247_n667_NOTT_99_n135(net238_c1,net238);
INTERCONNECT Split_255_n675_AND2T_89_n113(net239_c1,net239);
INTERCONNECT Split_263_n683_AND2T_57_n81(net240_c1,net240);
INTERCONNECT Split_271_n691_OR2T_30_n54(net241_c1,net241);
INTERCONNECT Split_319_n739_Split_320_n740(net242_c1,net242);
INTERCONNECT Split_327_n747_DFFT_137__FPB_n557(net243_c1,net243);
INTERCONNECT Split_248_n668_Split_249_n669(net244_c1,net244);
INTERCONNECT Split_256_n676_Split_257_n677(net245_c1,net245);
INTERCONNECT Split_264_n684_AND2T_19_n43(net246_c1,net246);
INTERCONNECT Split_272_n692_OR2T_33_n57(net247_c1,net247);
INTERCONNECT Split_328_n748_Split_329_n749(net248_c1,net248);
INTERCONNECT Split_249_n669_DFFT_154__FPB_n574(net249_c1,net249);
INTERCONNECT Split_257_n677_AND2T_15_n39(net250_c1,net250);
INTERCONNECT Split_265_n685_DFFT_136__FPB_n556(net251_c1,net251);
INTERCONNECT Split_273_n693_AND2T_38_n62(net252_c1,net252);
INTERCONNECT Split_329_n749_NOTT_16_n40(net253_c1,net253);
INTERCONNECT Split_258_n678_AND2T_62_n86(net254_c1,net254);
INTERCONNECT Split_266_n686_AND2T_22_n46(net255_c1,net255);
INTERCONNECT Split_274_n694_DFFT_194__FPB_n614(net256_c1,net256);
INTERCONNECT Split_259_n679_AND2T_42_n66(net257_c1,net257);
INTERCONNECT Split_267_n687_AND2T_25_n49(net258_c1,net258);
INTERCONNECT Split_275_n695_AND2T_89_n113(net259_c1,net259);
INTERCONNECT Split_268_n688_Split_269_n689(net260_c1,net260);
INTERCONNECT Split_276_n696_OR2T_60_n84(net261_c1,net261);
INTERCONNECT Split_269_n689_AND2T_28_n52(net262_c1,net262);
INTERCONNECT Split_277_n697_AND2T_65_n89(net263_c1,net263);
INTERCONNECT Split_278_n698_AND2T_43_n67(net264_c1,net264);
INTERCONNECT Split_279_n699_DFFT_170__FPB_n590(net265_c1,net265);
INTERCONNECT DFFT_106__PIPL_n154_DFFT_217__FPB_n637(net266_c1,net266);
INTERCONNECT DFFT_107__PIPL_n155_DFFT_225__FPB_n645(net267_c1,net267);
INTERCONNECT DFFT_108__PIPL_n156_DFFT_233__FPB_n653(net268_c1,net268);
INTERCONNECT DFFT_109__PIPL_n157_DFFT_240__FPB_n660(net269_c1,net269);
INTERCONNECT DFFT_110__FBL_n530_Split_316_n736(net270_c1,net270);
INTERCONNECT DFFT_111__FBL_n531_Split_317_n737(net271_c1,net271);
INTERCONNECT DFFT_120__FBL_n540_Split_325_n745(net272_c1,net272);
INTERCONNECT DFFT_112__FBL_n532_DFFT_187__FPB_n607(net273_c1,net273);
INTERCONNECT DFFT_121__FBL_n541_Split_328_n748(net274_c1,net274);
INTERCONNECT DFFT_113__FBL_n533_DFFT_191__FPB_n611(net275_c1,net275);
INTERCONNECT DFFT_114__FBL_n534_NOTT_100_n136(net276_c1,net276);
INTERCONNECT DFFT_115__FBL_n535_Split_HOLD_591(net277_c1,net277);
INTERCONNECT DFFT_116__FBL_n536_Split_318_n738(net278_c1,net278);
INTERCONNECT DFFT_117__FBL_n537_AND2T_103_n139(net279_c1,net279);
INTERCONNECT DFFT_118__FBL_n538_Split_319_n739(net280_c1,net280);
INTERCONNECT DFFT_119__FBL_n539_Split_322_n742(net281_c1,net281);
INTERCONNECT DFFT_104__FPB_n152_Split_310_n730(net282_c1,net282);
INTERCONNECT DFFT_105__FPB_n153_Split_313_n733(net283_c1,net283);
INTERCONNECT DFFT_180__FPB_n600_DFFT_181__FPB_n601(net284_c1,net284);
INTERCONNECT DFFT_181__FPB_n601_DFFT_182__FPB_n602(net285_c1,net285);
INTERCONNECT DFFT_182__FPB_n602_DFFT_183__FPB_n603(net286_c1,net286);
INTERCONNECT DFFT_190__FPB_n610_AND2T_75_n99(net287_c1,net287);
INTERCONNECT DFFT_191__FPB_n611_DFFT_192__FPB_n612(net288_c1,net288);
INTERCONNECT DFFT_183__FPB_n603_AND2T_70_n94(net289_c1,net289);
INTERCONNECT DFFT_200__FPB_n620_DFFT_201__FPB_n621(net290_c1,net290);
INTERCONNECT DFFT_192__FPB_n612_DFFT_193__FPB_n613(net291_c1,net291);
INTERCONNECT DFFT_184__FPB_n604_AND2T_71_n95(net292_c1,net292);
INTERCONNECT DFFT_201__FPB_n621_AND2T_83_n107(net293_c1,net293);
INTERCONNECT DFFT_193__FPB_n613_OR2T_76_n100(net294_c1,net294);
INTERCONNECT DFFT_185__FPB_n605_OR2T_73_n97(net295_c1,net295);
INTERCONNECT DFFT_210__FPB_n630_DFFT_211__FPB_n631(net296_c1,net296);
INTERCONNECT DFFT_202__FPB_n622_DFFT_203__FPB_n623(net297_c1,net297);
INTERCONNECT DFFT_122__FPB_n542_DFFT_112__FBL_n532(net298_c1,net298);
INTERCONNECT DFFT_194__FPB_n614_AND2T_79_n103(net299_c1,net299);
INTERCONNECT DFFT_186__FPB_n606_OR2T_74_n98(net300_c1,net300);
INTERCONNECT DFFT_130__FPB_n550_OR2T_23_n47(net301_c1,net301);
INTERCONNECT DFFT_211__FPB_n631_DFFT_212__FPB_n632(net302_c1,net302);
INTERCONNECT DFFT_203__FPB_n623_DFFT_204__FPB_n624(net303_c1,net303);
INTERCONNECT DFFT_187__FPB_n607_Split_HOLD_586(net304_c1,net304);
INTERCONNECT DFFT_123__FPB_n543_DFFT_113__FBL_n533(net305_c1,net305);
INTERCONNECT DFFT_195__FPB_n615_OR2T_82_n106(net306_c1,net306);
INTERCONNECT DFFT_131__FPB_n551_OR2T_24_n48(net307_c1,net307);
INTERCONNECT DFFT_220__FPB_n640_DFFT_221__FPB_n641(net308_c1,net308);
INTERCONNECT DFFT_212__FPB_n632_DFFT_213__FPB_n633(net309_c1,net309);
INTERCONNECT DFFT_196__FPB_n616_DFFT_197__FPB_n617(net310_c1,net310);
INTERCONNECT DFFT_188__FPB_n608_DFFT_189__FPB_n609(net311_c1,net311);
INTERCONNECT DFFT_132__FPB_n552_DFFT_133__FPB_n553(net312_c1,net312);
INTERCONNECT DFFT_124__FPB_n544_DFFT_116__FBL_n536(net313_c1,net313);
INTERCONNECT DFFT_204__FPB_n624_AND2T_84_n108(net314_c1,net314);
INTERCONNECT DFFT_140__FPB_n560_OR2T_30_n54(net315_c1,net315);
INTERCONNECT DFFT_221__FPB_n641_Split_HOLD_590(net316_c1,net316);
INTERCONNECT DFFT_213__FPB_n633_DFFT_214__FPB_n634(net317_c1,net317);
INTERCONNECT DFFT_197__FPB_n617_DFFT_198__FPB_n618(net318_c1,net318);
INTERCONNECT DFFT_189__FPB_n609_DFFT_190__FPB_n610(net319_c1,net319);
INTERCONNECT DFFT_133__FPB_n553_DFFT_134__FPB_n554(net320_c1,net320);
INTERCONNECT DFFT_125__FPB_n545_DFFT_117__FBL_n537(net321_c1,net321);
INTERCONNECT DFFT_205__FPB_n625_Split_HOLD_589(net322_c1,net322);
INTERCONNECT DFFT_141__FPB_n561_AND2T_32_n56(net323_c1,net323);
INTERCONNECT DFFT_230__FPB_n650_DFFT_231__FPB_n651(net324_c1,net324);
INTERCONNECT DFFT_222__FPB_n642_DFFT_223__FPB_n643(net325_c1,net325);
INTERCONNECT DFFT_214__FPB_n634_DFFT_215__FPB_n635(net326_c1,net326);
INTERCONNECT DFFT_198__FPB_n618_DFFT_199__FPB_n619(net327_c1,net327);
INTERCONNECT DFFT_142__FPB_n562_DFFT_143__FPB_n563(net328_c1,net328);
INTERCONNECT DFFT_134__FPB_n554_DFFT_135__FPB_n555(net329_c1,net329);
INTERCONNECT DFFT_126__FPB_n546_DFFT_120__FBL_n540(net330_c1,net330);
INTERCONNECT DFFT_206__FPB_n626_OR2T_90_n114(net331_c1,net331);
INTERCONNECT DFFT_150__FPB_n570_AND2T_44_n68(net332_c1,net332);
INTERCONNECT DFFT_231__FPB_n651_DFFT_232_state_obs1(net333_c1,net333);
INTERCONNECT DFFT_223__FPB_n643_DFFT_224_state_obs0(net334_c1,net334);
INTERCONNECT DFFT_207__FPB_n627_DFFT_208__FPB_n628(net335_c1,net335);
INTERCONNECT DFFT_199__FPB_n619_DFFT_200__FPB_n620(net336_c1,net336);
INTERCONNECT DFFT_127__FPB_n547_DFFT_121__FBL_n541(net337_c1,net337);
INTERCONNECT DFFT_215__FPB_n635_AND2T_94_n118(net338_c1,net338);
INTERCONNECT DFFT_151__FPB_n571_AND2T_45_n69(net339_c1,net339);
INTERCONNECT DFFT_143__FPB_n563_OR2T_33_n57(net340_c1,net340);
INTERCONNECT DFFT_135__FPB_n555_AND2T_25_n49(net341_c1,net341);
INTERCONNECT DFFT_240__FPB_n660_DFFT_241__FPB_n661(net342_c1,net342);
INTERCONNECT DFFT_216__FPB_n636_OR2T_96_n120(net343_c1,net343);
INTERCONNECT DFFT_208__FPB_n628_OR2T_92_n116(net344_c1,net344);
INTERCONNECT DFFT_160__FPB_n580_AND2T_53_n77(net345_c1,net345);
INTERCONNECT DFFT_152__FPB_n572_OR2T_50_n74(net346_c1,net346);
INTERCONNECT DFFT_144__FPB_n564_OR2T_35_n59(net347_c1,net347);
INTERCONNECT DFFT_136__FPB_n556_AND2T_26_n50(net348_c1,net348);
INTERCONNECT DFFT_128__FPB_n548_AND2T_14_n38(net349_c1,net349);
INTERCONNECT DFFT_241__FPB_n661_DFFT_242__FPB_n662(net350_c1,net350);
INTERCONNECT DFFT_233__FPB_n653_DFFT_234__FPB_n654(net351_c1,net351);
INTERCONNECT DFFT_225__FPB_n645_DFFT_226__FPB_n646(net352_c1,net352);
INTERCONNECT DFFT_217__FPB_n637_DFFT_218__FPB_n638(net353_c1,net353);
INTERCONNECT DFFT_209__FPB_n629_OR2T_93_n117(net354_c1,net354);
INTERCONNECT DFFT_161__FPB_n581_OR2T_55_n79(net355_c1,net355);
INTERCONNECT DFFT_153__FPB_n573_OR2T_52_n76(net356_c1,net356);
INTERCONNECT DFFT_145__FPB_n565_AND2T_36_n60(net357_c1,net357);
INTERCONNECT DFFT_137__FPB_n557_AND2T_27_n51(net358_c1,net358);
INTERCONNECT DFFT_129__FPB_n549_AND2T_18_n42(net359_c1,net359);
INTERCONNECT DFFT_242__FPB_n662_DFFT_243__FPB_n663(net360_c1,net360);
INTERCONNECT DFFT_234__FPB_n654_DFFT_235__FPB_n655(net361_c1,net361);
INTERCONNECT DFFT_226__FPB_n646_DFFT_227__FPB_n647(net362_c1,net362);
INTERCONNECT DFFT_218__FPB_n638_DFFT_219__FPB_n639(net363_c1,net363);
INTERCONNECT DFFT_162__FPB_n582_DFFT_163__FPB_n583(net364_c1,net364);
INTERCONNECT DFFT_154__FPB_n574_DFFT_155__FPB_n575(net365_c1,net365);
INTERCONNECT DFFT_138__FPB_n558_DFFT_139__FPB_n559(net366_c1,net366);
INTERCONNECT DFFT_170__FPB_n590_OR2T_60_n84(net367_c1,net367);
INTERCONNECT DFFT_146__FPB_n566_Split_HOLD_593(net368_c1,net368);
INTERCONNECT DFFT_243__FPB_n663_DFFT_244__FPB_n664(net369_c1,net369);
INTERCONNECT DFFT_235__FPB_n655_DFFT_236__FPB_n656(net370_c1,net370);
INTERCONNECT DFFT_227__FPB_n647_DFFT_228__FPB_n648(net371_c1,net371);
INTERCONNECT DFFT_219__FPB_n639_DFFT_220__FPB_n640(net372_c1,net372);
INTERCONNECT DFFT_171__FPB_n591_DFFT_172__FPB_n592(net373_c1,net373);
INTERCONNECT DFFT_163__FPB_n583_DFFT_164__FPB_n584(net374_c1,net374);
INTERCONNECT DFFT_155__FPB_n575_DFFT_156__FPB_n576(net375_c1,net375);
INTERCONNECT DFFT_139__FPB_n559_DFFT_140__FPB_n560(net376_c1,net376);
INTERCONNECT DFFT_147__FPB_n567_AND2T_39_n63(net377_c1,net377);
INTERCONNECT DFFT_244__FPB_n664_DFFT_245_state_obs3(net378_c1,net378);
INTERCONNECT DFFT_236__FPB_n656_DFFT_237__FPB_n657(net379_c1,net379);
INTERCONNECT DFFT_228__FPB_n648_DFFT_229__FPB_n649(net380_c1,net380);
INTERCONNECT DFFT_164__FPB_n584_DFFT_165__FPB_n585(net381_c1,net381);
INTERCONNECT DFFT_156__FPB_n576_DFFT_157__FPB_n577(net382_c1,net382);
INTERCONNECT DFFT_172__FPB_n592_AND2T_61_n85(net383_c1,net383);
INTERCONNECT DFFT_148__FPB_n568_AND2T_42_n66(net384_c1,net384);
INTERCONNECT DFFT_237__FPB_n657_DFFT_238__FPB_n658(net385_c1,net385);
INTERCONNECT DFFT_229__FPB_n649_DFFT_230__FPB_n650(net386_c1,net386);
INTERCONNECT DFFT_165__FPB_n585_DFFT_166__FPB_n586(net387_c1,net387);
INTERCONNECT DFFT_157__FPB_n577_DFFT_158__FPB_n578(net388_c1,net388);
INTERCONNECT DFFT_149__FPB_n569_DFFT_150__FPB_n570(net389_c1,net389);
INTERCONNECT DFFT_173__FPB_n593_AND2T_62_n86(net390_c1,net390);
INTERCONNECT DFFT_238__FPB_n658_DFFT_239_state_obs2(net391_c1,net391);
INTERCONNECT DFFT_158__FPB_n578_DFFT_159__FPB_n579(net392_c1,net392);
INTERCONNECT DFFT_174__FPB_n594_AND2T_64_n88(net393_c1,net393);
INTERCONNECT DFFT_166__FPB_n586_AND2T_56_n80(net394_c1,net394);
INTERCONNECT DFFT_167__FPB_n587_DFFT_168__FPB_n588(net395_c1,net395);
INTERCONNECT DFFT_159__FPB_n579_DFFT_160__FPB_n580(net396_c1,net396);
INTERCONNECT DFFT_175__FPB_n595_OR2T_66_n90(net397_c1,net397);
INTERCONNECT DFFT_168__FPB_n588_Split_HOLD_587(net398_c1,net398);
INTERCONNECT DFFT_176__FPB_n596_OR2T_68_n92(net399_c1,net399);
INTERCONNECT DFFT_177__FPB_n597_DFFT_178__FPB_n598(net400_c1,net400);
INTERCONNECT DFFT_169__FPB_n589_AND2T_59_n83(net401_c1,net401);
INTERCONNECT DFFT_178__FPB_n598_DFFT_179__FPB_n599(net402_c1,net402);
INTERCONNECT DFFT_179__FPB_n599_DFFT_180__FPB_n600(net403_c1,net403);
INTERCONNECT DFFT_224_state_obs0_state_obs0_Pad(net404_c1,state_obs0_Pad);
INTERCONNECT DFFT_232_state_obs1_state_obs1_Pad(net405_c1,state_obs1_Pad);
INTERCONNECT DFFT_239_state_obs2_state_obs2_Pad(net406_c1,state_obs2_Pad);
INTERCONNECT DFFT_245_state_obs3_state_obs3_Pad(net407_c1,state_obs3_Pad);
INTERCONNECT DFFT_97_state0_buf_DFFT_106__PIPL_n154(net408_c1,net408);
INTERCONNECT DFFT_98_state1_buf_DFFT_107__PIPL_n155(net409_c1,net409);
INTERCONNECT SplitCLK_0_493_SplitCLK_0_356(net410_c1,net410);
INTERCONNECT SplitCLK_0_493_SplitCLK_2_474(net411_c1,net411);
INTERCONNECT SplitCLK_2_492_DFFT_189__FPB_n609(net412_c1,net412);
INTERCONNECT SplitCLK_2_491_DFFT_158__FPB_n578(net413_c1,net413);
INTERCONNECT SplitCLK_2_490_DFFT_181__FPB_n601(net414_c1,net414);
INTERCONNECT SplitCLK_2_489_DFFT_148__FPB_n568(net415_c1,net415);
INTERCONNECT SplitCLK_4_488_DFFT_164__FPB_n584(net416_c1,net416);
INTERCONNECT SplitCLK_2_487_DFFT_155__FPB_n575(net417_c1,net417);
INTERCONNECT SplitCLK_4_486_DFFT_171__FPB_n591(net418_c1,net418);
INTERCONNECT SplitCLK_4_485_DFFT_162__FPB_n582(net419_c1,net419);
INTERCONNECT SplitCLK_2_484_DFFT_226__FPB_n646(net420_c1,net420);
INTERCONNECT SplitCLK_2_483_DFFT_131__FPB_n551(net421_c1,net421);
INTERCONNECT SplitCLK_2_482_DFFT_211__FPB_n631(net422_c1,net422);
INTERCONNECT SplitCLK_2_481_DFFT_121__FBL_n541(net423_c1,net423);
INTERCONNECT SplitCLK_4_480_DFFT_110__FBL_n530(net424_c1,net424);
INTERCONNECT SplitCLK_2_479_OR2T_48_n72(net425_c1,net425);
INTERCONNECT SplitCLK_2_478_AND2T_59_n83(net426_c1,net426);
INTERCONNECT SplitCLK_2_477_AND2T_26_n50(net427_c1,net427);
INTERCONNECT SplitCLK_2_476_AND2T_25_n49(net428_c1,net428);
INTERCONNECT SplitCLK_2_475_NOTT_8_n32(net429_c1,net429);
INTERCONNECT SplitCLK_2_474_SplitCLK_6_415(net430_c1,net430);
INTERCONNECT SplitCLK_2_474_SplitCLK_4_473(net431_c1,net431);
INTERCONNECT SplitCLK_4_473_SplitCLK_0_444(net432_c1,net432);
INTERCONNECT SplitCLK_4_473_SplitCLK_2_472(net433_c1,net433);
INTERCONNECT SplitCLK_2_472_SplitCLK_6_458(net434_c1,net434);
INTERCONNECT SplitCLK_2_472_SplitCLK_4_471(net435_c1,net435);
INTERCONNECT SplitCLK_4_471_SplitCLK_0_464(net436_c1,net436);
INTERCONNECT SplitCLK_4_471_SplitCLK_2_470(net437_c1,net437);
INTERCONNECT SplitCLK_2_470_SplitCLK_6_467(net438_c1,net438);
INTERCONNECT SplitCLK_2_470_SplitCLK_4_469(net439_c1,net439);
INTERCONNECT SplitCLK_4_469_SplitCLK_2_491(net440_c1,net440);
INTERCONNECT SplitCLK_4_469_SplitCLK_4_468(net441_c1,net441);
INTERCONNECT SplitCLK_4_468_DFFT_156__FPB_n576(net442_c1,net442);
INTERCONNECT SplitCLK_4_468_DFFT_157__FPB_n577(net443_c1,net443);
INTERCONNECT SplitCLK_6_467_SplitCLK_4_465(net444_c1,net444);
INTERCONNECT SplitCLK_6_467_SplitCLK_4_466(net445_c1,net445);
INTERCONNECT SplitCLK_4_466_DFFT_105__FPB_n153(net446_c1,net446);
INTERCONNECT SplitCLK_4_466_DFFT_159__FPB_n579(net447_c1,net447);
INTERCONNECT SplitCLK_4_465_DFFT_160__FPB_n580(net448_c1,net448);
INTERCONNECT SplitCLK_4_465_DFFT_183__FPB_n603(net449_c1,net449);
INTERCONNECT SplitCLK_0_464_SplitCLK_6_461(net450_c1,net450);
INTERCONNECT SplitCLK_0_464_SplitCLK_2_463(net451_c1,net451);
INTERCONNECT SplitCLK_2_463_SplitCLK_2_487(net452_c1,net452);
INTERCONNECT SplitCLK_2_463_SplitCLK_4_462(net453_c1,net453);
INTERCONNECT SplitCLK_4_462_DFFT_123__FPB_n543(net454_c1,net454);
INTERCONNECT SplitCLK_4_462_DFFT_182__FPB_n602(net455_c1,net455);
INTERCONNECT SplitCLK_6_461_SplitCLK_4_459(net456_c1,net456);
INTERCONNECT SplitCLK_6_461_SplitCLK_4_460(net457_c1,net457);
INTERCONNECT SplitCLK_4_460_DFFT_104__FPB_n152(net458_c1,net458);
INTERCONNECT SplitCLK_4_460_NOTT_99_n135(net459_c1,net459);
INTERCONNECT SplitCLK_4_459_DFFT_113__FBL_n533(net460_c1,net460);
INTERCONNECT SplitCLK_4_459_DFFT_163__FPB_n583(net461_c1,net461);
INTERCONNECT SplitCLK_6_458_SplitCLK_4_451(net462_c1,net462);
INTERCONNECT SplitCLK_6_458_SplitCLK_6_457(net463_c1,net463);
INTERCONNECT SplitCLK_6_457_SplitCLK_2_454(net464_c1,net464);
INTERCONNECT SplitCLK_6_457_SplitCLK_6_456(net465_c1,net465);
INTERCONNECT SplitCLK_6_456_SplitCLK_4_485(net466_c1,net466);
INTERCONNECT SplitCLK_6_456_SplitCLK_4_455(net467_c1,net467);
INTERCONNECT SplitCLK_4_455_AND2T_61_n85(net468_c1,net468);
INTERCONNECT SplitCLK_4_455_AND2T_53_n77(net469_c1,net469);
INTERCONNECT SplitCLK_2_454_SplitCLK_4_452(net470_c1,net470);
INTERCONNECT SplitCLK_2_454_SplitCLK_4_453(net471_c1,net471);
INTERCONNECT SplitCLK_4_453_OR2T_35_n59(net472_c1,net472);
INTERCONNECT SplitCLK_4_453_DFFT_172__FPB_n592(net473_c1,net473);
INTERCONNECT SplitCLK_4_452_OR2T_50_n74(net474_c1,net474);
INTERCONNECT SplitCLK_4_452_OR2T_51_n75(net475_c1,net475);
INTERCONNECT SplitCLK_4_451_SplitCLK_6_447(net476_c1,net476);
INTERCONNECT SplitCLK_4_451_SplitCLK_2_450(net477_c1,net477);
INTERCONNECT SplitCLK_2_450_SplitCLK_4_448(net478_c1,net478);
INTERCONNECT SplitCLK_2_450_SplitCLK_4_449(net479_c1,net479);
INTERCONNECT SplitCLK_4_449_NOTT_9_n33(net480_c1,net480);
INTERCONNECT SplitCLK_4_449_DFFT_149__FPB_n569(net481_c1,net481);
INTERCONNECT SplitCLK_4_448_AND2T_70_n94(net482_c1,net482);
INTERCONNECT SplitCLK_4_448_DFFT_166__FPB_n586(net483_c1,net483);
INTERCONNECT SplitCLK_6_447_SplitCLK_4_445(net484_c1,net484);
INTERCONNECT SplitCLK_6_447_SplitCLK_4_446(net485_c1,net485);
INTERCONNECT SplitCLK_4_446_OR2T_33_n57(net486_c1,net486);
INTERCONNECT SplitCLK_4_446_DFFT_142__FPB_n562(net487_c1,net487);
INTERCONNECT SplitCLK_4_445_AND2T_34_n58(net488_c1,net488);
INTERCONNECT SplitCLK_4_445_AND2T_44_n68(net489_c1,net489);
INTERCONNECT SplitCLK_0_444_SplitCLK_4_429(net490_c1,net490);
INTERCONNECT SplitCLK_0_444_SplitCLK_4_443(net491_c1,net491);
INTERCONNECT SplitCLK_4_443_SplitCLK_0_436(net492_c1,net492);
INTERCONNECT SplitCLK_4_443_SplitCLK_6_442(net493_c1,net493);
INTERCONNECT SplitCLK_6_442_SplitCLK_4_439(net494_c1,net494);
INTERCONNECT SplitCLK_6_442_SplitCLK_4_441(net495_c1,net495);
INTERCONNECT SplitCLK_4_441_SplitCLK_2_490(net496_c1,net496);
INTERCONNECT SplitCLK_4_441_SplitCLK_4_440(net497_c1,net497);
INTERCONNECT SplitCLK_4_440_DFFT_180__FPB_n600(net498_c1,net498);
INTERCONNECT SplitCLK_4_440_DFFT_179__FPB_n599(net499_c1,net499);
INTERCONNECT SplitCLK_4_439_SplitCLK_4_437(net500_c1,net500);
INTERCONNECT SplitCLK_4_439_SplitCLK_4_438(net501_c1,net501);
INTERCONNECT SplitCLK_4_438_DFFT_191__FPB_n611(net502_c1,net502);
INTERCONNECT SplitCLK_4_438_DFFT_192__FPB_n612(net503_c1,net503);
INTERCONNECT SplitCLK_4_437_DFFT_165__FPB_n585(net504_c1,net504);
INTERCONNECT SplitCLK_4_437_DFFT_193__FPB_n613(net505_c1,net505);
INTERCONNECT SplitCLK_0_436_SplitCLK_4_432(net506_c1,net506);
INTERCONNECT SplitCLK_0_436_SplitCLK_4_435(net507_c1,net507);
INTERCONNECT SplitCLK_4_435_SplitCLK_4_433(net508_c1,net508);
INTERCONNECT SplitCLK_4_435_SplitCLK_2_434(net509_c1,net509);
INTERCONNECT SplitCLK_2_434_OR2T_76_n100(net510_c1,net510);
INTERCONNECT SplitCLK_2_434_DFFT_178__FPB_n598(net511_c1,net511);
INTERCONNECT SplitCLK_4_433_DFFT_154__FPB_n574(net512_c1,net512);
INTERCONNECT SplitCLK_4_433_DFFT_177__FPB_n597(net513_c1,net513);
INTERCONNECT SplitCLK_4_432_SplitCLK_4_430(net514_c1,net514);
INTERCONNECT SplitCLK_4_432_SplitCLK_4_431(net515_c1,net515);
INTERCONNECT SplitCLK_4_431_AND2T_75_n99(net516_c1,net516);
INTERCONNECT SplitCLK_4_431_DFFT_167__FPB_n587(net517_c1,net517);
INTERCONNECT SplitCLK_4_430_DFFT_190__FPB_n610(net518_c1,net518);
INTERCONNECT SplitCLK_4_430_DFFT_168__FPB_n588(net519_c1,net519);
INTERCONNECT SplitCLK_4_429_SplitCLK_6_422(net520_c1,net520);
INTERCONNECT SplitCLK_4_429_SplitCLK_6_428(net521_c1,net521);
INTERCONNECT SplitCLK_6_428_SplitCLK_6_425(net522_c1,net522);
INTERCONNECT SplitCLK_6_428_SplitCLK_6_427(net523_c1,net523);
INTERCONNECT SplitCLK_6_427_SplitCLK_4_488(net524_c1,net524);
INTERCONNECT SplitCLK_6_427_SplitCLK_4_426(net525_c1,net525);
INTERCONNECT SplitCLK_4_426_AND2T_56_n80(net526_c1,net526);
INTERCONNECT SplitCLK_4_426_OR2T_69_n93(net527_c1,net527);
INTERCONNECT SplitCLK_6_425_SplitCLK_4_423(net528_c1,net528);
INTERCONNECT SplitCLK_6_425_SplitCLK_4_424(net529_c1,net529);
INTERCONNECT SplitCLK_4_424_DFFT_150__FPB_n570(net530_c1,net530);
INTERCONNECT SplitCLK_4_424_DFFT_143__FPB_n563(net531_c1,net531);
INTERCONNECT SplitCLK_4_423_OR2T_52_n76(net532_c1,net532);
INTERCONNECT SplitCLK_4_423_OR2T_54_n78(net533_c1,net533);
INTERCONNECT SplitCLK_6_422_SplitCLK_6_418(net534_c1,net534);
INTERCONNECT SplitCLK_6_422_SplitCLK_4_421(net535_c1,net535);
INTERCONNECT SplitCLK_4_421_SplitCLK_4_419(net536_c1,net536);
INTERCONNECT SplitCLK_4_421_SplitCLK_4_420(net537_c1,net537);
INTERCONNECT SplitCLK_4_420_OR2T_55_n79(net538_c1,net538);
INTERCONNECT SplitCLK_4_420_OR2T_68_n92(net539_c1,net539);
INTERCONNECT SplitCLK_4_419_DFFT_134__FPB_n554(net540_c1,net540);
INTERCONNECT SplitCLK_4_419_DFFT_135__FPB_n555(net541_c1,net541);
INTERCONNECT SplitCLK_6_418_SplitCLK_4_416(net542_c1,net542);
INTERCONNECT SplitCLK_6_418_SplitCLK_4_417(net543_c1,net543);
INTERCONNECT SplitCLK_4_417_OR2T_24_n48(net544_c1,net544);
INTERCONNECT SplitCLK_4_417_DFFT_161__FPB_n581(net545_c1,net545);
INTERCONNECT SplitCLK_4_416_OR2T_23_n47(net546_c1,net546);
INTERCONNECT SplitCLK_4_416_DFFT_153__FPB_n573(net547_c1,net547);
INTERCONNECT SplitCLK_6_415_SplitCLK_6_385(net548_c1,net548);
INTERCONNECT SplitCLK_6_415_SplitCLK_2_414(net549_c1,net549);
INTERCONNECT SplitCLK_2_414_SplitCLK_6_399(net550_c1,net550);
INTERCONNECT SplitCLK_2_414_SplitCLK_4_413(net551_c1,net551);
INTERCONNECT SplitCLK_4_413_SplitCLK_0_406(net552_c1,net552);
INTERCONNECT SplitCLK_4_413_SplitCLK_2_412(net553_c1,net553);
INTERCONNECT SplitCLK_2_412_SplitCLK_2_409(net554_c1,net554);
INTERCONNECT SplitCLK_2_412_SplitCLK_4_411(net555_c1,net555);
INTERCONNECT SplitCLK_4_411_SplitCLK_4_486(net556_c1,net556);
INTERCONNECT SplitCLK_4_411_SplitCLK_4_410(net557_c1,net557);
INTERCONNECT SplitCLK_4_410_AND2T_18_n42(net558_c1,net558);
INTERCONNECT SplitCLK_4_410_DFFT_129__FPB_n549(net559_c1,net559);
INTERCONNECT SplitCLK_2_409_SplitCLK_4_407(net560_c1,net560);
INTERCONNECT SplitCLK_2_409_SplitCLK_4_408(net561_c1,net561);
INTERCONNECT SplitCLK_4_408_DFFT_114__FBL_n534(net562_c1,net562);
INTERCONNECT SplitCLK_4_408_NOTT_100_n136(net563_c1,net563);
INTERCONNECT SplitCLK_4_407_DFFT_118__FBL_n538(net564_c1,net564);
INTERCONNECT SplitCLK_4_407_DFFT_119__FBL_n539(net565_c1,net565);
INTERCONNECT SplitCLK_0_406_SplitCLK_6_402(net566_c1,net566);
INTERCONNECT SplitCLK_0_406_SplitCLK_4_405(net567_c1,net567);
INTERCONNECT SplitCLK_4_405_SplitCLK_4_403(net568_c1,net568);
INTERCONNECT SplitCLK_4_405_SplitCLK_4_404(net569_c1,net569);
INTERCONNECT SplitCLK_4_404_DFFT_152__FPB_n572(net570_c1,net570);
INTERCONNECT SplitCLK_4_404_DFFT_144__FPB_n564(net571_c1,net571);
INTERCONNECT SplitCLK_4_403_AND2T_12_n36(net572_c1,net572);
INTERCONNECT SplitCLK_4_403_OR2T_49_n73(net573_c1,net573);
INTERCONNECT SplitCLK_6_402_SplitCLK_4_400(net574_c1,net574);
INTERCONNECT SplitCLK_6_402_SplitCLK_0_401(net575_c1,net575);
INTERCONNECT SplitCLK_0_401_AND2T_36_n60(net576_c1,net576);
INTERCONNECT SplitCLK_0_401_DFFT_174__FPB_n594(net577_c1,net577);
INTERCONNECT SplitCLK_4_400_AND2T_43_n67(net578_c1,net578);
INTERCONNECT SplitCLK_4_400_DFFT_146__FPB_n566(net579_c1,net579);
INTERCONNECT SplitCLK_6_399_SplitCLK_4_392(net580_c1,net580);
INTERCONNECT SplitCLK_6_399_SplitCLK_2_398(net581_c1,net581);
INTERCONNECT SplitCLK_2_398_SplitCLK_0_395(net582_c1,net582);
INTERCONNECT SplitCLK_2_398_SplitCLK_6_397(net583_c1,net583);
INTERCONNECT SplitCLK_6_397_SplitCLK_4_480(net584_c1,net584);
INTERCONNECT SplitCLK_6_397_SplitCLK_4_396(net585_c1,net585);
INTERCONNECT SplitCLK_4_396_DFFT_220__FPB_n640(net586_c1,net586);
INTERCONNECT SplitCLK_4_396_DFFT_219__FPB_n639(net587_c1,net587);
INTERCONNECT SplitCLK_0_395_SplitCLK_4_393(net588_c1,net588);
INTERCONNECT SplitCLK_0_395_SplitCLK_0_394(net589_c1,net589);
INTERCONNECT SplitCLK_0_394_DFFT_223__FPB_n643(net590_c1,net590);
INTERCONNECT SplitCLK_0_394_DFFT_224_state_obs0(net591_c1,net591);
INTERCONNECT SplitCLK_4_393_DFFT_221__FPB_n641(net592_c1,net592);
INTERCONNECT SplitCLK_4_393_DFFT_218__FPB_n638(net593_c1,net593);
INTERCONNECT SplitCLK_4_392_SplitCLK_0_388(net594_c1,net594);
INTERCONNECT SplitCLK_4_392_SplitCLK_4_391(net595_c1,net595);
INTERCONNECT SplitCLK_4_391_SplitCLK_4_389(net596_c1,net596);
INTERCONNECT SplitCLK_4_391_SplitCLK_4_390(net597_c1,net597);
INTERCONNECT SplitCLK_4_390_DFFT_97_state0_buf(net598_c1,net598);
INTERCONNECT SplitCLK_4_390_NOTT_101_n137(net599_c1,net599);
INTERCONNECT SplitCLK_4_389_DFFT_106__PIPL_n154(net600_c1,net600);
INTERCONNECT SplitCLK_4_389_DFFT_115__FBL_n535(net601_c1,net601);
INTERCONNECT SplitCLK_0_388_SplitCLK_4_386(net602_c1,net602);
INTERCONNECT SplitCLK_0_388_SplitCLK_0_387(net603_c1,net603);
INTERCONNECT SplitCLK_0_387_DFFT_222__FPB_n642(net604_c1,net604);
INTERCONNECT SplitCLK_0_387_DFFT_232_state_obs1(net605_c1,net605);
INTERCONNECT SplitCLK_4_386_DFFT_217__FPB_n637(net606_c1,net606);
INTERCONNECT SplitCLK_4_386_DFFT_229__FPB_n649(net607_c1,net607);
INTERCONNECT SplitCLK_6_385_SplitCLK_6_370(net608_c1,net608);
INTERCONNECT SplitCLK_6_385_SplitCLK_4_384(net609_c1,net609);
INTERCONNECT SplitCLK_4_384_SplitCLK_0_377(net610_c1,net610);
INTERCONNECT SplitCLK_4_384_SplitCLK_4_383(net611_c1,net611);
INTERCONNECT SplitCLK_4_383_SplitCLK_6_380(net612_c1,net612);
INTERCONNECT SplitCLK_4_383_SplitCLK_4_382(net613_c1,net613);
INTERCONNECT SplitCLK_4_382_SplitCLK_2_479(net614_c1,net614);
INTERCONNECT SplitCLK_4_382_SplitCLK_4_381(net615_c1,net615);
INTERCONNECT SplitCLK_4_381_AND2T_15_n39(net616_c1,net616);
INTERCONNECT SplitCLK_4_381_AND2T_45_n69(net617_c1,net617);
INTERCONNECT SplitCLK_6_380_SplitCLK_4_378(net618_c1,net618);
INTERCONNECT SplitCLK_6_380_SplitCLK_0_379(net619_c1,net619);
INTERCONNECT SplitCLK_0_379_AND2T_38_n62(net620_c1,net620);
INTERCONNECT SplitCLK_0_379_DFFT_170__FPB_n590(net621_c1,net621);
INTERCONNECT SplitCLK_4_378_OR2T_41_n65(net622_c1,net622);
INTERCONNECT SplitCLK_4_378_OR2T_60_n84(net623_c1,net623);
INTERCONNECT SplitCLK_0_377_SplitCLK_6_373(net624_c1,net624);
INTERCONNECT SplitCLK_0_377_SplitCLK_4_376(net625_c1,net625);
INTERCONNECT SplitCLK_4_376_SplitCLK_4_374(net626_c1,net626);
INTERCONNECT SplitCLK_4_376_SplitCLK_4_375(net627_c1,net627);
INTERCONNECT SplitCLK_4_375_AND2T_57_n81(net628_c1,net628);
INTERCONNECT SplitCLK_4_375_OR2T_67_n91(net629_c1,net629);
INTERCONNECT SplitCLK_4_374_AND2T_31_n55(net630_c1,net630);
INTERCONNECT SplitCLK_4_374_AND2T_28_n52(net631_c1,net631);
INTERCONNECT SplitCLK_6_373_SplitCLK_4_371(net632_c1,net632);
INTERCONNECT SplitCLK_6_373_SplitCLK_4_372(net633_c1,net633);
INTERCONNECT SplitCLK_4_372_AND2T_37_n61(net634_c1,net634);
INTERCONNECT SplitCLK_4_372_OR2T_66_n90(net635_c1,net635);
INTERCONNECT SplitCLK_4_371_AND2T_40_n64(net636_c1,net636);
INTERCONNECT SplitCLK_4_371_AND2T_47_n71(net637_c1,net637);
INTERCONNECT SplitCLK_6_370_SplitCLK_0_363(net638_c1,net638);
INTERCONNECT SplitCLK_6_370_SplitCLK_6_369(net639_c1,net639);
INTERCONNECT SplitCLK_6_369_SplitCLK_6_366(net640_c1,net640);
INTERCONNECT SplitCLK_6_369_SplitCLK_6_368(net641_c1,net641);
INTERCONNECT SplitCLK_6_368_SplitCLK_2_484(net642_c1,net642);
INTERCONNECT SplitCLK_6_368_SplitCLK_4_367(net643_c1,net643);
INTERCONNECT SplitCLK_4_367_AND2T_64_n88(net644_c1,net644);
INTERCONNECT SplitCLK_4_367_DFFT_175__FPB_n595(net645_c1,net645);
INTERCONNECT SplitCLK_6_366_SplitCLK_4_364(net646_c1,net646);
INTERCONNECT SplitCLK_6_366_SplitCLK_4_365(net647_c1,net647);
INTERCONNECT SplitCLK_4_365_DFFT_230__FPB_n650(net648_c1,net648);
INTERCONNECT SplitCLK_4_365_DFFT_227__FPB_n647(net649_c1,net649);
INTERCONNECT SplitCLK_4_364_DFFT_231__FPB_n651(net650_c1,net650);
INTERCONNECT SplitCLK_4_364_DFFT_228__FPB_n648(net651_c1,net651);
INTERCONNECT SplitCLK_0_363_SplitCLK_6_359(net652_c1,net652);
INTERCONNECT SplitCLK_0_363_SplitCLK_4_362(net653_c1,net653);
INTERCONNECT SplitCLK_4_362_SplitCLK_4_360(net654_c1,net654);
INTERCONNECT SplitCLK_4_362_SplitCLK_4_361(net655_c1,net655);
INTERCONNECT SplitCLK_4_361_AND2T_65_n89(net656_c1,net656);
INTERCONNECT SplitCLK_4_361_DFFT_225__FPB_n645(net657_c1,net657);
INTERCONNECT SplitCLK_4_360_DFFT_111__FBL_n531(net658_c1,net658);
INTERCONNECT SplitCLK_4_360_DFFT_128__FPB_n548(net659_c1,net659);
INTERCONNECT SplitCLK_6_359_SplitCLK_4_357(net660_c1,net660);
INTERCONNECT SplitCLK_6_359_SplitCLK_0_358(net661_c1,net661);
INTERCONNECT SplitCLK_0_358_DFFT_239_state_obs2(net662_c1,net662);
INTERCONNECT SplitCLK_0_358_DFFT_237__FPB_n657(net663_c1,net663);
INTERCONNECT SplitCLK_4_357_DFFT_107__PIPL_n155(net664_c1,net664);
INTERCONNECT SplitCLK_4_357_DFFT_238__FPB_n658(net665_c1,net665);
INTERCONNECT SplitCLK_0_356_SplitCLK_6_297(net666_c1,net666);
INTERCONNECT SplitCLK_0_356_SplitCLK_4_355(net667_c1,net667);
INTERCONNECT SplitCLK_4_355_SplitCLK_0_326(net668_c1,net668);
INTERCONNECT SplitCLK_4_355_SplitCLK_2_354(net669_c1,net669);
INTERCONNECT SplitCLK_2_354_SplitCLK_6_340(net670_c1,net670);
INTERCONNECT SplitCLK_2_354_SplitCLK_4_353(net671_c1,net671);
INTERCONNECT SplitCLK_4_353_SplitCLK_4_346(net672_c1,net672);
INTERCONNECT SplitCLK_4_353_SplitCLK_2_352(net673_c1,net673);
INTERCONNECT SplitCLK_2_352_SplitCLK_6_349(net674_c1,net674);
INTERCONNECT SplitCLK_2_352_SplitCLK_4_351(net675_c1,net675);
INTERCONNECT SplitCLK_4_351_SplitCLK_2_492(net676_c1,net676);
INTERCONNECT SplitCLK_4_351_SplitCLK_4_350(net677_c1,net677);
INTERCONNECT SplitCLK_4_350_DFFT_212__FPB_n632(net678_c1,net678);
INTERCONNECT SplitCLK_4_350_DFFT_213__FPB_n633(net679_c1,net679);
INTERCONNECT SplitCLK_6_349_SplitCLK_4_347(net680_c1,net680);
INTERCONNECT SplitCLK_6_349_SplitCLK_0_348(net681_c1,net681);
INTERCONNECT SplitCLK_0_348_DFFT_169__FPB_n589(net682_c1,net682);
INTERCONNECT SplitCLK_0_348_DFFT_188__FPB_n608(net683_c1,net683);
INTERCONNECT SplitCLK_4_347_AND2T_77_n101(net684_c1,net684);
INTERCONNECT SplitCLK_4_347_DFFT_187__FPB_n607(net685_c1,net685);
INTERCONNECT SplitCLK_4_346_SplitCLK_0_343(net686_c1,net686);
INTERCONNECT SplitCLK_4_346_SplitCLK_2_345(net687_c1,net687);
INTERCONNECT SplitCLK_2_345_SplitCLK_2_482(net688_c1,net688);
INTERCONNECT SplitCLK_2_345_SplitCLK_4_344(net689_c1,net689);
INTERCONNECT SplitCLK_4_344_DFFT_210__FPB_n630(net690_c1,net690);
INTERCONNECT SplitCLK_4_344_DFFT_214__FPB_n634(net691_c1,net691);
INTERCONNECT SplitCLK_0_343_SplitCLK_4_341(net692_c1,net692);
INTERCONNECT SplitCLK_0_343_SplitCLK_0_342(net693_c1,net693);
INTERCONNECT SplitCLK_0_342_AND2T_94_n118(net694_c1,net694);
INTERCONNECT SplitCLK_0_342_OR2T_82_n106(net695_c1,net695);
INTERCONNECT SplitCLK_4_341_DFFT_112__FBL_n532(net696_c1,net696);
INTERCONNECT SplitCLK_4_341_DFFT_215__FPB_n635(net697_c1,net697);
INTERCONNECT SplitCLK_6_340_SplitCLK_0_333(net698_c1,net698);
INTERCONNECT SplitCLK_6_340_SplitCLK_6_339(net699_c1,net699);
INTERCONNECT SplitCLK_6_339_SplitCLK_6_336(net700_c1,net700);
INTERCONNECT SplitCLK_6_339_SplitCLK_2_338(net701_c1,net701);
INTERCONNECT SplitCLK_2_338_SplitCLK_2_476(net702_c1,net702);
INTERCONNECT SplitCLK_2_338_SplitCLK_4_337(net703_c1,net703);
INTERCONNECT SplitCLK_4_337_DFFT_132__FPB_n552(net704_c1,net704);
INTERCONNECT SplitCLK_4_337_DFFT_133__FPB_n553(net705_c1,net705);
INTERCONNECT SplitCLK_6_336_SplitCLK_4_334(net706_c1,net706);
INTERCONNECT SplitCLK_6_336_SplitCLK_4_335(net707_c1,net707);
INTERCONNECT SplitCLK_4_335_OR2T_30_n54(net708_c1,net708);
INTERCONNECT SplitCLK_4_335_DFFT_130__FPB_n550(net709_c1,net709);
INTERCONNECT SplitCLK_4_334_DFFT_140__FPB_n560(net710_c1,net710);
INTERCONNECT SplitCLK_4_334_OR2T_81_n105(net711_c1,net711);
INTERCONNECT SplitCLK_0_333_SplitCLK_4_329(net712_c1,net712);
INTERCONNECT SplitCLK_0_333_SplitCLK_4_332(net713_c1,net713);
INTERCONNECT SplitCLK_4_332_SplitCLK_4_330(net714_c1,net714);
INTERCONNECT SplitCLK_4_332_SplitCLK_4_331(net715_c1,net715);
INTERCONNECT SplitCLK_4_331_DFFT_138__FPB_n558(net716_c1,net716);
INTERCONNECT SplitCLK_4_331_DFFT_139__FPB_n559(net717_c1,net717);
INTERCONNECT SplitCLK_4_330_OR2T_93_n117(net718_c1,net718);
INTERCONNECT SplitCLK_4_330_DFFT_176__FPB_n596(net719_c1,net719);
INTERCONNECT SplitCLK_4_329_SplitCLK_4_327(net720_c1,net720);
INTERCONNECT SplitCLK_4_329_SplitCLK_4_328(net721_c1,net721);
INTERCONNECT SplitCLK_4_328_DFFT_141__FPB_n561(net722_c1,net722);
INTERCONNECT SplitCLK_4_328_DFFT_195__FPB_n615(net723_c1,net723);
INTERCONNECT SplitCLK_4_327_AND2T_22_n46(net724_c1,net724);
INTERCONNECT SplitCLK_4_327_AND2T_85_n109(net725_c1,net725);
INTERCONNECT SplitCLK_0_326_SplitCLK_6_311(net726_c1,net726);
INTERCONNECT SplitCLK_0_326_SplitCLK_4_325(net727_c1,net727);
INTERCONNECT SplitCLK_4_325_SplitCLK_4_318(net728_c1,net728);
INTERCONNECT SplitCLK_4_325_SplitCLK_2_324(net729_c1,net729);
INTERCONNECT SplitCLK_2_324_SplitCLK_6_321(net730_c1,net730);
INTERCONNECT SplitCLK_2_324_SplitCLK_4_323(net731_c1,net731);
INTERCONNECT SplitCLK_4_323_SplitCLK_2_475(net732_c1,net732);
INTERCONNECT SplitCLK_4_323_SplitCLK_4_322(net733_c1,net733);
INTERCONNECT SplitCLK_4_322_DFFT_196__FPB_n616(net734_c1,net734);
INTERCONNECT SplitCLK_4_322_DFFT_197__FPB_n617(net735_c1,net735);
INTERCONNECT SplitCLK_6_321_SplitCLK_4_319(net736_c1,net736);
INTERCONNECT SplitCLK_6_321_SplitCLK_0_320(net737_c1,net737);
INTERCONNECT SplitCLK_0_320_DFFT_122__FPB_n542(net738_c1,net738);
INTERCONNECT SplitCLK_0_320_DFFT_209__FPB_n629(net739_c1,net739);
INTERCONNECT SplitCLK_4_319_DFFT_124__FPB_n544(net740_c1,net740);
INTERCONNECT SplitCLK_4_319_DFFT_127__FPB_n547(net741_c1,net741);
INTERCONNECT SplitCLK_4_318_SplitCLK_0_314(net742_c1,net742);
INTERCONNECT SplitCLK_4_318_SplitCLK_6_317(net743_c1,net743);
INTERCONNECT SplitCLK_6_317_SplitCLK_4_315(net744_c1,net744);
INTERCONNECT SplitCLK_6_317_SplitCLK_4_316(net745_c1,net745);
INTERCONNECT SplitCLK_4_316_AND2T_83_n107(net746_c1,net746);
INTERCONNECT SplitCLK_4_316_DFFT_198__FPB_n618(net747_c1,net747);
INTERCONNECT SplitCLK_4_315_DFFT_199__FPB_n619(net748_c1,net748);
INTERCONNECT SplitCLK_4_315_DFFT_201__FPB_n621(net749_c1,net749);
INTERCONNECT SplitCLK_0_314_SplitCLK_4_312(net750_c1,net750);
INTERCONNECT SplitCLK_0_314_SplitCLK_0_313(net751_c1,net751);
INTERCONNECT SplitCLK_0_313_DFFT_116__FBL_n536(net752_c1,net752);
INTERCONNECT SplitCLK_0_313_DFFT_126__FPB_n546(net753_c1,net753);
INTERCONNECT SplitCLK_4_312_DFFT_200__FPB_n620(net754_c1,net754);
INTERCONNECT SplitCLK_4_312_DFFT_125__FPB_n545(net755_c1,net755);
INTERCONNECT SplitCLK_6_311_SplitCLK_4_304(net756_c1,net756);
INTERCONNECT SplitCLK_6_311_SplitCLK_4_310(net757_c1,net757);
INTERCONNECT SplitCLK_4_310_SplitCLK_6_307(net758_c1,net758);
INTERCONNECT SplitCLK_4_310_SplitCLK_6_309(net759_c1,net759);
INTERCONNECT SplitCLK_6_309_SplitCLK_2_478(net760_c1,net760);
INTERCONNECT SplitCLK_6_309_SplitCLK_4_308(net761_c1,net761);
INTERCONNECT SplitCLK_4_308_AND2T_84_n108(net762_c1,net762);
INTERCONNECT SplitCLK_4_308_DFFT_204__FPB_n624(net763_c1,net763);
INTERCONNECT SplitCLK_6_307_SplitCLK_4_305(net764_c1,net764);
INTERCONNECT SplitCLK_6_307_SplitCLK_4_306(net765_c1,net765);
INTERCONNECT SplitCLK_4_306_OR2T_92_n116(net766_c1,net766);
INTERCONNECT SplitCLK_4_306_DFFT_208__FPB_n628(net767_c1,net767);
INTERCONNECT SplitCLK_4_305_AND2T_71_n95(net768_c1,net768);
INTERCONNECT SplitCLK_4_305_DFFT_207__FPB_n627(net769_c1,net769);
INTERCONNECT SplitCLK_4_304_SplitCLK_0_300(net770_c1,net770);
INTERCONNECT SplitCLK_4_304_SplitCLK_4_303(net771_c1,net771);
INTERCONNECT SplitCLK_4_303_SplitCLK_4_301(net772_c1,net772);
INTERCONNECT SplitCLK_4_303_SplitCLK_4_302(net773_c1,net773);
INTERCONNECT SplitCLK_4_302_AND2T_86_n110(net774_c1,net774);
INTERCONNECT SplitCLK_4_302_DFFT_203__FPB_n623(net775_c1,net775);
INTERCONNECT SplitCLK_4_301_DFFT_202__FPB_n622(net776_c1,net776);
INTERCONNECT SplitCLK_4_301_DFFT_117__FBL_n537(net777_c1,net777);
INTERCONNECT SplitCLK_0_300_SplitCLK_4_298(net778_c1,net778);
INTERCONNECT SplitCLK_0_300_SplitCLK_0_299(net779_c1,net779);
INTERCONNECT SplitCLK_0_299_OR2T_74_n98(net780_c1,net780);
INTERCONNECT SplitCLK_0_299_DFFT_186__FPB_n606(net781_c1,net781);
INTERCONNECT SplitCLK_4_298_AND2T_103_n139(net782_c1,net782);
INTERCONNECT SplitCLK_4_298_DFFT_184__FPB_n604(net783_c1,net783);
INTERCONNECT SplitCLK_6_297_SplitCLK_0_267(net784_c1,net784);
INTERCONNECT SplitCLK_6_297_SplitCLK_2_296(net785_c1,net785);
INTERCONNECT SplitCLK_2_296_SplitCLK_6_281(net786_c1,net786);
INTERCONNECT SplitCLK_2_296_SplitCLK_4_295(net787_c1,net787);
INTERCONNECT SplitCLK_4_295_SplitCLK_0_288(net788_c1,net788);
INTERCONNECT SplitCLK_4_295_SplitCLK_4_294(net789_c1,net789);
INTERCONNECT SplitCLK_4_294_SplitCLK_6_291(net790_c1,net790);
INTERCONNECT SplitCLK_4_294_SplitCLK_4_293(net791_c1,net791);
INTERCONNECT SplitCLK_4_293_SplitCLK_2_483(net792_c1,net792);
INTERCONNECT SplitCLK_4_293_SplitCLK_4_292(net793_c1,net793);
INTERCONNECT SplitCLK_4_292_AND2T_19_n43(net794_c1,net794);
INTERCONNECT SplitCLK_4_292_OR2T_58_n82(net795_c1,net795);
INTERCONNECT SplitCLK_6_291_SplitCLK_4_289(net796_c1,net796);
INTERCONNECT SplitCLK_6_291_SplitCLK_4_290(net797_c1,net797);
INTERCONNECT SplitCLK_4_290_AND2T_46_n70(net798_c1,net798);
INTERCONNECT SplitCLK_4_290_AND2T_39_n63(net799_c1,net799);
INTERCONNECT SplitCLK_4_289_OR2T_80_n104(net800_c1,net800);
INTERCONNECT SplitCLK_4_289_DFFT_147__FPB_n567(net801_c1,net801);
INTERCONNECT SplitCLK_0_288_SplitCLK_4_284(net802_c1,net802);
INTERCONNECT SplitCLK_0_288_SplitCLK_4_287(net803_c1,net803);
INTERCONNECT SplitCLK_4_287_SplitCLK_4_285(net804_c1,net804);
INTERCONNECT SplitCLK_4_287_SplitCLK_4_286(net805_c1,net805);
INTERCONNECT SplitCLK_4_286_AND2T_32_n56(net806_c1,net806);
INTERCONNECT SplitCLK_4_286_AND2T_79_n103(net807_c1,net807);
INTERCONNECT SplitCLK_4_285_OR2T_29_n53(net808_c1,net808);
INTERCONNECT SplitCLK_4_285_AND2T_78_n102(net809_c1,net809);
INTERCONNECT SplitCLK_4_284_SplitCLK_0_282(net810_c1,net810);
INTERCONNECT SplitCLK_4_284_SplitCLK_4_283(net811_c1,net811);
INTERCONNECT SplitCLK_4_283_AND2T_20_n44(net812_c1,net812);
INTERCONNECT SplitCLK_4_283_NOTT_11_n35(net813_c1,net813);
INTERCONNECT SplitCLK_0_282_AND2T_14_n38(net814_c1,net814);
INTERCONNECT SplitCLK_0_282_DFFT_194__FPB_n614(net815_c1,net815);
INTERCONNECT SplitCLK_6_281_SplitCLK_4_274(net816_c1,net816);
INTERCONNECT SplitCLK_6_281_SplitCLK_6_280(net817_c1,net817);
INTERCONNECT SplitCLK_6_280_SplitCLK_6_277(net818_c1,net818);
INTERCONNECT SplitCLK_6_280_SplitCLK_2_279(net819_c1,net819);
INTERCONNECT SplitCLK_2_279_SplitCLK_2_489(net820_c1,net820);
INTERCONNECT SplitCLK_2_279_SplitCLK_4_278(net821_c1,net821);
INTERCONNECT SplitCLK_4_278_AND2T_42_n66(net822_c1,net822);
INTERCONNECT SplitCLK_4_278_AND2T_62_n86(net823_c1,net823);
INTERCONNECT SplitCLK_6_277_SplitCLK_4_275(net824_c1,net824);
INTERCONNECT SplitCLK_6_277_SplitCLK_4_276(net825_c1,net825);
INTERCONNECT SplitCLK_4_276_DFFT_245_state_obs3(net826_c1,net826);
INTERCONNECT SplitCLK_4_276_DFFT_98_state1_buf(net827_c1,net827);
INTERCONNECT SplitCLK_4_275_DFFT_108__PIPL_n156(net828_c1,net828);
INTERCONNECT SplitCLK_4_275_DFFT_233__FPB_n653(net829_c1,net829);
INTERCONNECT SplitCLK_4_274_SplitCLK_6_270(net830_c1,net830);
INTERCONNECT SplitCLK_4_274_SplitCLK_4_273(net831_c1,net831);
INTERCONNECT SplitCLK_4_273_SplitCLK_4_271(net832_c1,net832);
INTERCONNECT SplitCLK_4_273_SplitCLK_4_272(net833_c1,net833);
INTERCONNECT SplitCLK_4_272_AND2T_89_n113(net834_c1,net834);
INTERCONNECT SplitCLK_4_272_DFFT_173__FPB_n593(net835_c1,net835);
INTERCONNECT SplitCLK_4_271_DFFT_206__FPB_n626(net836_c1,net836);
INTERCONNECT SplitCLK_4_271_DFFT_145__FPB_n565(net837_c1,net837);
INTERCONNECT SplitCLK_6_270_SplitCLK_4_268(net838_c1,net838);
INTERCONNECT SplitCLK_6_270_SplitCLK_4_269(net839_c1,net839);
INTERCONNECT SplitCLK_4_269_DFFT_234__FPB_n654(net840_c1,net840);
INTERCONNECT SplitCLK_4_269_NOTT_95_n119(net841_c1,net841);
INTERCONNECT SplitCLK_4_268_NOTT_16_n40(net842_c1,net842);
INTERCONNECT SplitCLK_4_268_DFFT_235__FPB_n655(net843_c1,net843);
INTERCONNECT SplitCLK_0_267_SplitCLK_6_252(net844_c1,net844);
INTERCONNECT SplitCLK_0_267_SplitCLK_4_266(net845_c1,net845);
INTERCONNECT SplitCLK_4_266_SplitCLK_0_259(net846_c1,net846);
INTERCONNECT SplitCLK_4_266_SplitCLK_2_265(net847_c1,net847);
INTERCONNECT SplitCLK_2_265_SplitCLK_6_262(net848_c1,net848);
INTERCONNECT SplitCLK_2_265_SplitCLK_2_264(net849_c1,net849);
INTERCONNECT SplitCLK_2_264_SplitCLK_2_477(net850_c1,net850);
INTERCONNECT SplitCLK_2_264_SplitCLK_4_263(net851_c1,net851);
INTERCONNECT SplitCLK_4_263_AND2T_72_n96(net852_c1,net852);
INTERCONNECT SplitCLK_4_263_DFFT_136__FPB_n556(net853_c1,net853);
INTERCONNECT SplitCLK_6_262_SplitCLK_4_260(net854_c1,net854);
INTERCONNECT SplitCLK_6_262_SplitCLK_4_261(net855_c1,net855);
INTERCONNECT SplitCLK_4_261_AND2T_17_n41(net856_c1,net856);
INTERCONNECT SplitCLK_4_261_NOTT_10_n34(net857_c1,net857);
INTERCONNECT SplitCLK_4_260_OR2T_73_n97(net858_c1,net858);
INTERCONNECT SplitCLK_4_260_DFFT_185__FPB_n605(net859_c1,net859);
INTERCONNECT SplitCLK_0_259_SplitCLK_6_255(net860_c1,net860);
INTERCONNECT SplitCLK_0_259_SplitCLK_4_258(net861_c1,net861);
INTERCONNECT SplitCLK_4_258_SplitCLK_4_256(net862_c1,net862);
INTERCONNECT SplitCLK_4_258_SplitCLK_4_257(net863_c1,net863);
INTERCONNECT SplitCLK_4_257_DFFT_151__FPB_n571(net864_c1,net864);
INTERCONNECT SplitCLK_4_257_OR2T_88_n112(net865_c1,net865);
INTERCONNECT SplitCLK_4_256_DFFT_205__FPB_n625(net866_c1,net866);
INTERCONNECT SplitCLK_4_256_NOTT_102_n138(net867_c1,net867);
INTERCONNECT SplitCLK_6_255_SplitCLK_4_253(net868_c1,net868);
INTERCONNECT SplitCLK_6_255_SplitCLK_4_254(net869_c1,net869);
INTERCONNECT SplitCLK_4_254_AND2T_27_n51(net870_c1,net870);
INTERCONNECT SplitCLK_4_254_OR2T_91_n115(net871_c1,net871);
INTERCONNECT SplitCLK_4_253_AND2T_87_n111(net872_c1,net872);
INTERCONNECT SplitCLK_4_253_OR2T_90_n114(net873_c1,net873);
INTERCONNECT SplitCLK_6_252_SplitCLK_4_245(net874_c1,net874);
INTERCONNECT SplitCLK_6_252_SplitCLK_2_251(net875_c1,net875);
INTERCONNECT SplitCLK_2_251_SplitCLK_6_248(net876_c1,net876);
INTERCONNECT SplitCLK_2_251_SplitCLK_2_250(net877_c1,net877);
INTERCONNECT SplitCLK_2_250_SplitCLK_2_481(net878_c1,net878);
INTERCONNECT SplitCLK_2_250_SplitCLK_4_249(net879_c1,net879);
INTERCONNECT SplitCLK_4_249_AND2T_63_n87(net880_c1,net880);
INTERCONNECT SplitCLK_4_249_DFFT_137__FPB_n557(net881_c1,net881);
INTERCONNECT SplitCLK_6_248_SplitCLK_4_246(net882_c1,net882);
INTERCONNECT SplitCLK_6_248_SplitCLK_4_247(net883_c1,net883);
INTERCONNECT SplitCLK_4_247_NOTT_13_n37(net884_c1,net884);
INTERCONNECT SplitCLK_4_247_DFFT_236__FPB_n656(net885_c1,net885);
INTERCONNECT SplitCLK_4_246_DFFT_240__FPB_n660(net886_c1,net886);
INTERCONNECT SplitCLK_4_246_OR2T_96_n120(net887_c1,net887);
INTERCONNECT SplitCLK_4_245_SplitCLK_6_241(net888_c1,net888);
INTERCONNECT SplitCLK_4_245_SplitCLK_2_244(net889_c1,net889);
INTERCONNECT SplitCLK_2_244_SplitCLK_4_242(net890_c1,net890);
INTERCONNECT SplitCLK_2_244_SplitCLK_0_243(net891_c1,net891);
INTERCONNECT SplitCLK_0_243_DFFT_109__PIPL_n157(net892_c1,net892);
INTERCONNECT SplitCLK_0_243_DFFT_216__FPB_n636(net893_c1,net893);
INTERCONNECT SplitCLK_4_242_AND2T_21_n45(net894_c1,net894);
INTERCONNECT SplitCLK_4_242_DFFT_120__FBL_n540(net895_c1,net895);
INTERCONNECT SplitCLK_6_241_SplitCLK_4_239(net896_c1,net896);
INTERCONNECT SplitCLK_6_241_SplitCLK_4_240(net897_c1,net897);
INTERCONNECT SplitCLK_4_240_DFFT_241__FPB_n661(net898_c1,net898);
INTERCONNECT SplitCLK_4_240_DFFT_242__FPB_n662(net899_c1,net899);
INTERCONNECT SplitCLK_4_239_DFFT_243__FPB_n663(net900_c1,net900);
INTERCONNECT SplitCLK_4_239_DFFT_244__FPB_n664(net901_c1,net901);
INTERCONNECT GCLK_Pad_SplitCLK_0_493(GCLK_Pad,net902);
INTERCONNECT Split_HOLD_586_DFFT_188__FPB_n608(net903_c1,net903);
INTERCONNECT Split_HOLD_587_DFFT_169__FPB_n589(net904_c1,net904);
INTERCONNECT Split_HOLD_588_AND2T_87_n111(net905_c1,net905);
INTERCONNECT Split_HOLD_589_AND2T_87_n111(net906_c1,net906);
INTERCONNECT Split_HOLD_590_DFFT_222__FPB_n642(net907_c1,net907);
INTERCONNECT Split_HOLD_591_NOTT_101_n137(net908_c1,net908);
INTERCONNECT Split_HOLD_592_DFFT_216__FPB_n636(net909_c1,net909);
INTERCONNECT Split_HOLD_593_AND2T_38_n62(net910_c1,net910);

endmodule
