module TAP_route(
input GCLK_Pad,
input TMS_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output state_obs2_Pad,
output state_obs3_Pad);

wire TMS_Pad;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire TRST_Pad;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire state_obs0_Pad;
wire net383_c1;
wire state_obs1_Pad;
wire net384_c1;
wire state_obs2_Pad;
wire net385_c1;
wire state_obs3_Pad;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire net486_c1;
wire net486;
wire net487_c1;
wire net487;
wire net488_c1;
wire net488;
wire net489_c1;
wire net489;
wire net490_c1;
wire net490;
wire net491_c1;
wire net491;
wire net492_c1;
wire net492;
wire net493_c1;
wire net493;
wire net494_c1;
wire net494;
wire net495_c1;
wire net495;
wire net496_c1;
wire net496;
wire net497_c1;
wire net497;
wire net498_c1;
wire net498;
wire net499_c1;
wire net499;
wire net500_c1;
wire net500;
wire net501_c1;
wire net501;
wire net502_c1;
wire net502;
wire net503_c1;
wire net503;
wire net504_c1;
wire net504;
wire net505_c1;
wire net505;
wire net506_c1;
wire net506;
wire net507_c1;
wire net507;
wire net508_c1;
wire net508;
wire net509_c1;
wire net509;
wire net510_c1;
wire net510;
wire net511_c1;
wire net511;
wire net512_c1;
wire net512;
wire net513_c1;
wire net513;
wire net514_c1;
wire net514;
wire net515_c1;
wire net515;
wire net516_c1;
wire net516;
wire net517_c1;
wire net517;
wire net518_c1;
wire net518;
wire net519_c1;
wire net519;
wire net520_c1;
wire net520;
wire net521_c1;
wire net521;
wire net522_c1;
wire net522;
wire net523_c1;
wire net523;
wire net524_c1;
wire net524;
wire net525_c1;
wire net525;
wire net526_c1;
wire net526;
wire net527_c1;
wire net527;
wire net528_c1;
wire net528;
wire net529_c1;
wire net529;
wire net530_c1;
wire net530;
wire net531_c1;
wire net531;
wire net532_c1;
wire net532;
wire net533_c1;
wire net533;
wire net534_c1;
wire net534;
wire net535_c1;
wire net535;
wire net536_c1;
wire net536;
wire net537_c1;
wire net537;
wire net538_c1;
wire net538;
wire net539_c1;
wire net539;
wire net540_c1;
wire net540;
wire net541_c1;
wire net541;
wire net542_c1;
wire net542;
wire net543_c1;
wire net543;
wire net544_c1;
wire net544;
wire net545_c1;
wire net545;
wire net546_c1;
wire net546;
wire net547_c1;
wire net547;
wire net548_c1;
wire net548;
wire net549_c1;
wire net549;
wire net550_c1;
wire net550;
wire net551_c1;
wire net551;
wire net552_c1;
wire net552;
wire net553_c1;
wire net553;
wire net554_c1;
wire net554;
wire net555_c1;
wire net555;
wire net556_c1;
wire net556;
wire net557_c1;
wire net557;
wire net558_c1;
wire net558;
wire net559_c1;
wire net559;
wire net560_c1;
wire net560;
wire net561_c1;
wire net561;
wire net562_c1;
wire net562;
wire net563_c1;
wire net563;
wire net564_c1;
wire net564;
wire net565_c1;
wire net565;
wire net566_c1;
wire net566;
wire net567_c1;
wire net567;
wire net568_c1;
wire net568;
wire net569_c1;
wire net569;
wire net570_c1;
wire net570;
wire net571_c1;
wire net571;
wire net572_c1;
wire net572;
wire net573_c1;
wire net573;
wire net574_c1;
wire net574;
wire net575_c1;
wire net575;
wire net576_c1;
wire net576;
wire net577_c1;
wire net577;
wire net578_c1;
wire net578;
wire net579_c1;
wire net579;
wire net580_c1;
wire net580;
wire net581_c1;
wire net581;
wire net582_c1;
wire net582;
wire net583_c1;
wire net583;
wire net584_c1;
wire net584;
wire net585_c1;
wire net585;
wire net586_c1;
wire net586;
wire net587_c1;
wire net587;
wire net588_c1;
wire net588;
wire net589_c1;
wire net589;
wire net590_c1;
wire net590;
wire net591_c1;
wire net591;
wire net592_c1;
wire net592;
wire net593_c1;
wire net593;
wire net594_c1;
wire net594;
wire net595_c1;
wire net595;
wire net596_c1;
wire net596;
wire net597_c1;
wire net597;
wire net598_c1;
wire net598;
wire net599_c1;
wire net599;
wire net600_c1;
wire net600;
wire net601_c1;
wire net601;
wire net602_c1;
wire net602;
wire net603_c1;
wire net603;
wire net604_c1;
wire net604;
wire net605_c1;
wire net605;
wire net606_c1;
wire net606;
wire net607_c1;
wire net607;
wire net608_c1;
wire net608;
wire net609_c1;
wire net609;
wire net610_c1;
wire net610;
wire net611_c1;
wire net611;
wire net612_c1;
wire net612;
wire net613_c1;
wire net613;
wire net614_c1;
wire net614;
wire net615_c1;
wire net615;
wire net616_c1;
wire net616;
wire net617_c1;
wire net617;
wire net618_c1;
wire net618;
wire net619_c1;
wire net619;
wire net620_c1;
wire net620;
wire net621_c1;
wire net621;
wire net622_c1;
wire net622;
wire net623_c1;
wire net623;
wire net624_c1;
wire net624;
wire net625_c1;
wire net625;
wire net626_c1;
wire net626;
wire net627_c1;
wire net627;
wire net628_c1;
wire net628;
wire net629_c1;
wire net629;
wire net630_c1;
wire net630;
wire net631_c1;
wire net631;
wire net632_c1;
wire net632;
wire net633_c1;
wire net633;
wire net634_c1;
wire net634;
wire net635_c1;
wire net635;
wire net636_c1;
wire net636;
wire net637_c1;
wire net637;
wire net638_c1;
wire net638;
wire net639_c1;
wire net639;
wire net640_c1;
wire net640;
wire net641_c1;
wire net641;
wire net642_c1;
wire net642;
wire net643_c1;
wire net643;
wire net644_c1;
wire net644;
wire net645_c1;
wire net645;
wire net646_c1;
wire net646;
wire net647_c1;
wire net647;
wire net648_c1;
wire net648;
wire net649_c1;
wire net649;
wire net650_c1;
wire net650;
wire net651_c1;
wire net651;
wire net652_c1;
wire net652;
wire net653_c1;
wire net653;
wire net654_c1;
wire net654;
wire net655_c1;
wire net655;
wire net656_c1;
wire net656;
wire net657_c1;
wire net657;
wire net658_c1;
wire net658;
wire net659_c1;
wire net659;
wire net660_c1;
wire net660;
wire net661_c1;
wire net661;
wire net662_c1;
wire net662;
wire net663_c1;
wire net663;
wire net664_c1;
wire net664;
wire net665_c1;
wire net665;
wire net666_c1;
wire net666;
wire net667_c1;
wire net667;
wire net668_c1;
wire net668;
wire net669_c1;
wire net669;
wire net670_c1;
wire net670;
wire net671_c1;
wire net671;
wire net672_c1;
wire net672;
wire net673_c1;
wire net673;
wire net674_c1;
wire net674;
wire net675_c1;
wire net675;
wire net676_c1;
wire net676;
wire net677_c1;
wire net677;
wire net678_c1;
wire net678;
wire net679_c1;
wire net679;
wire net680_c1;
wire net680;
wire net681_c1;
wire net681;
wire net682_c1;
wire net682;
wire net683_c1;
wire net683;
wire net684_c1;
wire net684;
wire net685_c1;
wire net685;
wire net686_c1;
wire net686;
wire net687_c1;
wire net687;
wire net688_c1;
wire net688;
wire net689_c1;
wire net689;
wire net690_c1;
wire net690;
wire net691_c1;
wire net691;
wire net692_c1;
wire net692;
wire net693_c1;
wire net693;
wire net694_c1;
wire net694;
wire net695_c1;
wire net695;
wire net696_c1;
wire net696;
wire net697_c1;
wire net697;
wire net698_c1;
wire net698;
wire net699_c1;
wire net699;
wire net700_c1;
wire net700;
wire net701_c1;
wire net701;
wire net702_c1;
wire net702;
wire net703_c1;
wire net703;
wire net704_c1;
wire net704;
wire net705_c1;
wire net705;
wire net706_c1;
wire net706;
wire net707_c1;
wire net707;
wire net708_c1;
wire net708;
wire net709_c1;
wire net709;
wire net710_c1;
wire net710;
wire net711_c1;
wire net711;
wire net712_c1;
wire net712;
wire net713_c1;
wire net713;
wire net714_c1;
wire net714;
wire net715_c1;
wire net715;
wire net716_c1;
wire net716;
wire net717_c1;
wire net717;
wire net718_c1;
wire net718;
wire net719_c1;
wire net719;
wire net720_c1;
wire net720;
wire net721_c1;
wire net721;
wire net722_c1;
wire net722;
wire net723_c1;
wire net723;
wire net724_c1;
wire net724;
wire net725_c1;
wire net725;
wire net726_c1;
wire net726;
wire net727_c1;
wire net727;
wire net728_c1;
wire net728;
wire net729_c1;
wire net729;
wire net730_c1;
wire net730;
wire net731_c1;
wire net731;
wire net732_c1;
wire net732;
wire net733_c1;
wire net733;
wire net734_c1;
wire net734;
wire net735_c1;
wire net735;
wire net736_c1;
wire net736;
wire net737_c1;
wire net737;
wire net738_c1;
wire net738;
wire net739_c1;
wire net739;
wire net740_c1;
wire net740;
wire net741_c1;
wire net741;
wire net742_c1;
wire net742;
wire net743_c1;
wire net743;
wire net744_c1;
wire net744;
wire net745_c1;
wire net745;
wire net746_c1;
wire net746;
wire net747_c1;
wire net747;
wire net748_c1;
wire net748;
wire net749_c1;
wire net749;
wire net750_c1;
wire net750;
wire net751_c1;
wire net751;
wire net752_c1;
wire net752;
wire net753_c1;
wire net753;
wire net754_c1;
wire net754;
wire net755_c1;
wire net755;
wire net756_c1;
wire net756;
wire net757_c1;
wire net757;
wire net758_c1;
wire net758;
wire net759_c1;
wire net759;
wire net760_c1;
wire net760;
wire net761_c1;
wire net761;
wire net762_c1;
wire net762;
wire net763_c1;
wire net763;
wire net764_c1;
wire net764;
wire net765_c1;
wire net765;
wire net766_c1;
wire net766;
wire net767_c1;
wire net767;
wire net768_c1;
wire net768;
wire net769_c1;
wire net769;
wire net770_c1;
wire net770;
wire net771_c1;
wire net771;
wire net772_c1;
wire net772;
wire net773_c1;
wire net773;
wire net774_c1;
wire net774;
wire net775_c1;
wire net775;
wire net776_c1;
wire net776;
wire net777_c1;
wire net777;
wire net778_c1;
wire net778;
wire net779_c1;
wire net779;
wire net780_c1;
wire net780;
wire net781_c1;
wire net781;
wire net782_c1;
wire net782;
wire net783_c1;
wire net783;
wire net784_c1;
wire net784;
wire net785_c1;
wire net785;
wire net786_c1;
wire net786;
wire net787_c1;
wire net787;
wire net788_c1;
wire net788;
wire net789_c1;
wire net789;
wire net790_c1;
wire net790;
wire net791_c1;
wire net791;
wire net792_c1;
wire net792;
wire net793_c1;
wire net793;
wire net794_c1;
wire net794;
wire net795_c1;
wire net795;
wire net796_c1;
wire net796;
wire net797_c1;
wire net797;
wire net798_c1;
wire net798;
wire net799_c1;
wire net799;
wire net800_c1;
wire net800;
wire net801_c1;
wire net801;
wire net802_c1;
wire net802;
wire net803_c1;
wire net803;
wire net804_c1;
wire net804;
wire net805_c1;
wire net805;
wire net806_c1;
wire net806;
wire net807_c1;
wire net807;
wire net808_c1;
wire net808;
wire net809_c1;
wire net809;
wire net810_c1;
wire net810;
wire net811_c1;
wire net811;
wire net812_c1;
wire net812;
wire net813_c1;
wire net813;
wire net814_c1;
wire net814;
wire net815_c1;
wire net815;
wire net816_c1;
wire net816;
wire net817_c1;
wire net817;
wire net818_c1;
wire net818;
wire net819_c1;
wire net819;
wire net820_c1;
wire net820;
wire net821_c1;
wire net821;
wire net822_c1;
wire net822;
wire net823_c1;
wire net823;
wire net824_c1;
wire net824;
wire net825_c1;
wire net825;
wire net826_c1;
wire net826;
wire net827_c1;
wire net827;
wire net828_c1;
wire net828;
wire net829_c1;
wire net829;
wire net830_c1;
wire net830;
wire net831_c1;
wire net831;
wire net832_c1;
wire net832;
wire net833_c1;
wire net833;
wire net834_c1;
wire net834;
wire net835_c1;
wire net835;
wire net836_c1;
wire net836;
wire net837_c1;
wire net837;
wire net838_c1;
wire net838;
wire net839_c1;
wire net839;
wire net840_c1;
wire net840;
wire net841_c1;
wire net841;
wire net842_c1;
wire net842;
wire net843_c1;
wire net843;
wire net844_c1;
wire net844;
wire net845_c1;
wire net845;
wire net846_c1;
wire net846;
wire net847_c1;
wire net847;
wire net848_c1;
wire net848;
wire net849_c1;
wire net849;
wire net850_c1;
wire net850;
wire net851_c1;
wire net851;
wire net852_c1;
wire net852;
wire net853_c1;
wire net853;
wire net854_c1;
wire net854;
wire net855_c1;
wire net855;
wire net856_c1;
wire net856;
wire net857_c1;
wire net857;
wire net858_c1;
wire net858;
wire net859_c1;
wire net859;
wire net860_c1;
wire net860;
wire net861_c1;
wire net861;
wire GCLK_Pad;
wire net862;
wire net863_c1;
wire net863;
wire net864_c1;
wire net864;
wire net865_c1;
wire net865;
wire net866_c1;
wire net866;
wire net867_c1;
wire net867;
wire net868_c1;
wire net868;

DFFT DFFT_99__FPB_n135(net658,net173,net267_c1);
DFFT DFFT_199__FPB_n589(net724,net378,net380_c1);
DFFT DFFT_209_state_obs0(net572,net381,net382_c1);
XOR2T XOR2T_48_n72(net634,net142,net285,net30_c1);
DFFT DFFT_229_state_obs3(net806,net332,net385_c1);
DFFT DFFT_100__PIPL_n136(net574,net4,net254_c1);
NOTT NOTT_8_n32(net546,net250,net2_c1);
NOTT NOTT_9_n33(net421,net178,net4_c1);
DFFT DFFT_101__PIPL_n137(net586,net10,net255_c1);
DFFT DFFT_102__PIPL_n138(net807,net18,net256_c1);
AND2T AND2T_20_n44(net766,net191,net132,net13_c1);
AND2T AND2T_21_n45(net558,net160,net170,net17_c1);
AND2T AND2T_30_n54(net780,net100,net297,net21_c1);
AND2T AND2T_22_n46(net788,net204,net234,net22_c1);
AND2T AND2T_14_n38(net794,net249,net172,net23_c1);
AND2T AND2T_31_n55(net420,net112,net239,net26_c1);
AND2T AND2T_15_n39(net800,net137,net291,net28_c1);
AND2T AND2T_40_n64(net542,net180,net302,net31_c1);
AND2T AND2T_32_n56(net822,net106,net303,net32_c1);
AND2T AND2T_24_n48(net789,net182,net223,net33_c1);
AND2T AND2T_41_n65(net762,net193,net159,net36_c1);
AND2T AND2T_25_n49(net419,net190,net304,net38_c1);
AND2T AND2T_26_n50(net778,net201,net188,net5_c1);
AND2T AND2T_42_n66(net474,net206,net317,net42_c1);
AND2T AND2T_19_n43(net600,net107,net97,net9_c1);
AND2T AND2T_43_n67(net418,net226,net324,net47_c1);
AND2T AND2T_35_n59(net560,net195,net192,net48_c1);
AND2T AND2T_36_n60(net614,net122,net279,net11_c1);
AND2T AND2T_60_n84(net668,net224,net352,net50_c1);
AND2T AND2T_44_n68(net763,net47,net217,net52_c1);
AND2T AND2T_29_n53(net470,net210,net290,net16_c1);
AND2T AND2T_61_n85(net774,net125,net184,net54_c1);
AND2T AND2T_53_n77(net417,net51,net294,net55_c1);
AND2T AND2T_45_n69(net596,net117,net331,net56_c1);
AND2T AND2T_70_n94(net690,net243,net335,net57_c1);
AND2T AND2T_62_n86(net828,net229,net310,net58_c1);
AND2T AND2T_47_n71(net608,net109,net30,net24_c1);
AND2T AND2T_39_n63(net476,net20,net43,net25_c1);
AND2T AND2T_71_n95(net696,net57,net199,net60_c1);
AND2T AND2T_63_n87(net834,net116,net316,net61_c1);
AND2T AND2T_56_n80(net416,net62,net337,net29_c1);
AND2T AND2T_57_n81(net415,net197,net110,net34_c1);
AND2T AND2T_58_n82(net775,net205,net242,net40_c1);
AND2T AND2T_74_n98(net816,net151,net342,net67_c1);
AND2T AND2T_69_n93(net492,net49,net329,net53_c1);
DFFT DFFT_103__PIPL_n139(net848,net1,net257_c1);
OR2T OR2T_16_n40(net767,net213,net298,net1_c1);
OR2T OR2T_33_n57(net781,net32,net26,net37_c1);
OR2T OR2T_50_n74(net464,net35,net295,net41_c1);
OR2T OR2T_34_n58(net528,net214,net275,net43_c1);
OR2T OR2T_27_n51(net768,net5,net269,net8_c1);
OR2T OR2T_51_n75(net462,net41,net25,net46_c1);
OR2T OR2T_28_n52(net612,net8,net271,net12_c1);
OR2T OR2T_52_n76(net465,net46,net301,net51_c1);
OR2T OR2T_37_n61(net477,net219,net289,net15_c1);
OR2T OR2T_46_n70(net414,net215,net211,net19_c1);
OR2T OR2T_38_n62(net554,net15,net296,net20_c1);
OR2T OR2T_54_n78(net518,net134,net141,net59_c1);
OR2T OR2T_55_n79(net529,net131,net300,net62_c1);
OR2T OR2T_72_n96(net738,net60,net202,net63_c1);
OR2T OR2T_64_n88(net530,net130,net126,net64_c1);
OR2T OR2T_49_n73(net609,net19,net288,net35_c1);
OR2T OR2T_73_n97(net748,net63,net136,net65_c1);
OR2T OR2T_65_n89(net682,net64,net323,net66_c1);
OR2T OR2T_66_n90(net413,net66,net330,net39_c1);
OR2T OR2T_67_n91(net659,net39,net336,net44_c1);
OR2T OR2T_59_n83(net817,net40,net34,net45_c1);
OR2T OR2T_75_n99(net412,net67,net220,net68_c1);
OR2T OR2T_68_n92(net502,net44,net29,net49_c1);
NOTT NOTT_10_n34(net561,net241,net7_c1);
NOTT NOTT_11_n35(net411,net186,net10_c1);
NOTT NOTT_12_n36(net547,net253,net14_c1);
NOTT NOTT_13_n37(net410,net218,net18_c1);
NOTT NOTT_23_n47(net409,net168,net27_c1);
NOTT NOTT_17_n41(net664,net108,net3_c1);
NOTT NOTT_18_n42(net531,net232,net6_c1);
AND2T AND2T_82_n106(net694,net80,net356,net84_c1);
AND2T AND2T_83_n107(net712,net146,net370,net87_c1);
AND2T AND2T_76_n100(net736,net203,net351,net69_c1);
AND2T AND2T_92_n116(net725,net86,net354,net88_c1);
AND2T AND2T_84_n108(net732,net129,net376,net89_c1);
AND2T AND2T_77_n101(net842,net21,net357,net70_c1);
AND2T AND2T_93_n120(net601,net233,net174,net75_c1);
AND2T AND2T_85_n109(net408,net121,net350,net90_c1);
AND2T AND2T_86_n110(net832,net73,net355,net71_c1);
AND2T AND2T_78_n102(net407,net212,net362,net72_c1);
AND2T AND2T_94_n121(net548,net14,net360,net78_c1);
AND2T AND2T_96_n123(net406,net209,net364,net85_c1);
DFFT DFFT_110__FBL_n500(net854,net278,net258_c1);
DFFT DFFT_111__FBL_n501(net568,net284,net259_c1);
DFFT DFFT_104__FBL_n494(net405,net55,net260_c1);
DFFT DFFT_120__FPB_n510(net769,net22,net269_c1);
DFFT DFFT_112__FPB_n502(net622,net221,net268_c1);
DFFT DFFT_200__FPB_n590(net718,net380,net354_c1);
DFFT DFFT_105__FBL_n495(net678,net207,net261_c1);
DFFT DFFT_121__FPB_n511(net615,net13,net271_c1);
DFFT DFFT_113__FPB_n503(net855,net225,net270_c1);
DFFT DFFT_201__FPB_n591(net559,net150,net360_c1);
DFFT DFFT_106__FBL_n496(net580,net268,net262_c1);
DFFT DFFT_210__FPB_n600(net623,net255,net272_c1);
DFFT DFFT_130__FPB_n520(net524,net315,net275_c1);
DFFT DFFT_122__FPB_n512(net450,net147,net273_c1);
DFFT DFFT_114__FPB_n504(net635,net139,net274_c1);
DFFT DFFT_202__FPB_n592(net581,net262,net364_c1);
DFFT DFFT_107__FBL_n497(net404,net270,net263_c1);
DFFT DFFT_211__FPB_n601(net628,net272,net276_c1);
DFFT DFFT_131__FPB_n521(net613,net238,net279_c1);
DFFT DFFT_123__FPB_n513(net458,net868,net277_c1);
DFFT DFFT_115__FPB_n505(net860,net145,net278_c1);
DFFT DFFT_203__FPB_n593(net573,net254,net367_c1);
DFFT DFFT_108__FBL_n498(net512,net124,net264_c1);
DFFT DFFT_220__FPB_n610(net804,net326,net280_c1);
DFFT DFFT_212__FPB_n602(net626,net276,net281_c1);
DFFT DFFT_140__FPB_n530(net843,net169,net285_c1);
DFFT DFFT_132__FPB_n522(net516,net152,net282_c1);
DFFT DFFT_124__FPB_n514(net403,net277,net283_c1);
DFFT DFFT_116__FPB_n506(net402,net216,net284_c1);
DFFT DFFT_204__FPB_n594(net569,net867,net371_c1);
DFFT DFFT_109__FBL_n499(net640,net274,net265_c1);
DFFT DFFT_221__FPB_n611(net795,net280,net286_c1);
DFFT DFFT_213__FPB_n603(net629,net281,net287_c1);
DFFT DFFT_141__FPB_n531(net401,net24,net288_c1);
DFFT DFFT_133__FPB_n523(net517,net282,net289_c1);
DFFT DFFT_125__FPB_n515(net459,net866,net290_c1);
DFFT DFFT_117__FPB_n507(net801,net251,net291_c1);
DFFT DFFT_205__FPB_n595(net587,net371,net374_c1);
DFFT DFFT_222__FPB_n612(net792,net286,net292_c1);
DFFT DFFT_214__FPB_n604(net638,net864,net293_c1);
DFFT DFFT_150__FPB_n540(net438,net341,net294_c1);
DFFT DFFT_142__FPB_n532(net475,net42,net295_c1);
DFFT DFFT_134__FPB_n524(net555,net48,net296_c1);
DFFT DFFT_126__FPB_n516(net779,net92,net297_c1);
DFFT DFFT_118__FPB_n508(net602,net156,net298_c1);
DFFT DFFT_206__FPB_n596(net584,net374,net377_c1);
DFFT DFFT_215__FPB_n605(net639,net293,net299_c1);
DFFT DFFT_151__FPB_n541(net519,net140,net300_c1);
DFFT DFFT_143__FPB_n533(net400,net16,net301_c1);
DFFT DFFT_135__FPB_n525(net543,net244,net302_c1);
DFFT DFFT_127__FPB_n517(net835,net127,net303_c1);
DFFT DFFT_119__FPB_n509(net549,net248,net304_c1);
DFFT DFFT_207__FPB_n597(net585,net377,net379_c1);
OR2T OR2T_80_n104(net697,net74,net68,net77_c1);
OR2T OR2T_81_n105(net695,net77,net366,net80_c1);
OR2T OR2T_90_n114(net744,net79,net361,net83_c1);
OR2T OR2T_91_n115(net722,net83,net365,net86_c1);
DFFT DFFT_224__FPB_n614(net858,net257,net305_c1);
DFFT DFFT_160__FPB_n550(net829,net135,net310_c1);
DFFT DFFT_152__FPB_n542(net439,net155,net306_c1);
DFFT DFFT_144__FPB_n534(net444,net179,net307_c1);
DFFT DFFT_136__FPB_n526(net399,net236,net308_c1);
DFFT DFFT_128__FPB_n518(net398,net231,net309_c1);
OR2T OR2T_87_n111(net597,net111,net99,net73_c1);
OR2T OR2T_79_n103(net737,net72,net69,net74_c1);
DFFT DFFT_208__FPB_n598(net575,net379,net381_c1);
OR2T OR2T_88_n112(net749,net71,net90,net76_c1);
OR2T OR2T_89_n113(net750,net76,net198,net79_c1);
DFFT DFFT_225__FPB_n615(net859,net305,net311_c1);
DFFT DFFT_217__FPB_n607(net397,net256,net312_c1);
DFFT DFFT_161__FPB_n551(net820,net194,net316_c1);
DFFT DFFT_153__FPB_n543(net448,net306,net313_c1);
DFFT DFFT_145__FPB_n535(net445,net307,net314_c1);
DFFT DFFT_137__FPB_n527(net471,net863,net317_c1);
DFFT DFFT_129__FPB_n519(net525,net309,net315_c1);
DFFT DFFT_226__FPB_n616(net861,net311,net318_c1);
DFFT DFFT_218__FPB_n608(net846,net312,net319_c1);
DFFT DFFT_170__FPB_n560(net490,net359,net320_c1);
DFFT DFFT_162__FPB_n552(net684,net119,net323_c1);
DFFT DFFT_154__FPB_n544(net451,net313,net321_c1);
DFFT DFFT_146__FPB_n536(net396,net314,net322_c1);
DFFT DFFT_138__FPB_n528(net463,net161,net324_c1);
DFFT DFFT_227__FPB_n617(net849,net318,net325_c1);
DFFT DFFT_219__FPB_n609(net805,net319,net326_c1);
DFFT DFFT_171__FPB_n561(net503,net320,net329_c1);
DFFT DFFT_163__FPB_n553(net683,net115,net330_c1);
DFFT DFFT_155__FPB_n545(net513,net321,net327_c1);
DFFT DFFT_147__FPB_n537(net434,net322,net328_c1);
DFFT DFFT_139__FPB_n529(net603,net158,net331_c1);
DFFT DFFT_228__FPB_n618(net847,net325,net332_c1);
DFFT DFFT_180__FPB_n570(net654,net369,net333_c1);
DFFT DFFT_172__FPB_n562(net679,net228,net335_c1);
DFFT DFFT_164__FPB_n554(net669,net50,net336_c1);
DFFT DFFT_156__FPB_n546(net491,net327,net337_c1);
DFFT DFFT_148__FPB_n538(net395,net328,net334_c1);
DFFT DFFT_181__FPB_n571(net498,net333,net338_c1);
DFFT DFFT_173__FPB_n563(net821,net163,net342_c1);
DFFT DFFT_165__FPB_n555(net486,net96,net339_c1);
DFFT DFFT_157__FPB_n547(net504,net149,net340_c1);
DFFT DFFT_149__FPB_n539(net435,net334,net341_c1);
DFFT DFFT_190__FPB_n580(net691,net144,net343_c1);
DFFT DFFT_182__FPB_n572(net655,net338,net344_c1);
DFFT DFFT_174__FPB_n564(net394,net162,net345_c1);
DFFT DFFT_166__FPB_n556(net487,net339,net346_c1);
DFFT DFFT_158__FPB_n548(net505,net340,net347_c1);
SPLITT Split_300_n690(net261,net144_c1,net228_c1);
SPLITT Split_301_n691(net263,net150_c1,net233_c1);
SPLITT Split_230_n620(net0,net91_c1,net173_c1);
SPLITT Split_310_n700(net171,net92_c1,net174_c1);
SPLITT Split_302_n692(net264,net153_c1,net237_c1);
SPLITT Split_231_n621(net91,net93_c1,net175_c1);
SPLITT Split_303_n693(net237,net160_c1,net241_c1);
SPLITT Split_232_n622(net2,net95_c1,net176_c1);
SPLITT Split_240_n630(net3,net94_c1,net177_c1);
SPLITT Split_304_n694(net153,net161_c1,net244_c1);
SPLITT Split_233_n623(net176,net97_c1,net178_c1);
SPLITT Split_241_n631(net177,net96_c1,net179_c1);
SPLITT Split_305_n695(net258,net164_c1,net247_c1);
SPLITT Split_234_n624(net95,net99_c1,net180_c1);
SPLITT Split_242_n632(net94,net98_c1,net181_c1);
SPLITT Split_250_n640(net128,net100_c1,net182_c1);
SPLITT Split_306_n696(net247,net168_c1,net249_c1);
SPLITT Split_235_n625(net7,net102_c1,net183_c1);
SPLITT Split_243_n633(net6,net103_c1,net184_c1);
SPLITT Split_251_n641(net33,net101_c1,net185_c1);
SPLITT Split_307_n697(net164,net169_c1,net251_c1);
SPLITT Split_236_n626(net183,net107_c1,net186_c1);
SPLITT Split_244_n634(net9,net105_c1,net187_c1);
SPLITT Split_252_n642(net185,net106_c1,net188_c1);
SPLITT Split_260_n650(net31,net104_c1,net189_c1);
SPLITT Split_308_n698(net259,net171_c1,net252_c1);
SPLITT Split_237_n627(net102,net111_c1,net190_c1);
SPLITT Split_245_n635(net187,net112_c1,net191_c1);
SPLITT Split_253_n643(net101,net110_c1,net192_c1);
SPLITT Split_261_n651(net189,net109_c1,net193_c1);
SPLITT Split_309_n699(net252,net172_c1,net253_c1);
SPLITT Split_238_n628(net23,net114_c1,net194_c1);
SPLITT Split_246_n636(net105,net117_c1,net195_c1);
SPLITT Split_254_n644(net38,net113_c1,net196_c1);
SPLITT Split_262_n652(net104,net116_c1,net197_c1);
SPLITT Split_270_n660(net58,net115_c1,net198_c1);
SPLITT Split_239_n629(net28,net121_c1,net199_c1);
SPLITT Split_247_n637(net17,net118_c1,net200_c1);
SPLITT Split_255_n645(net196,net122_c1,net201_c1);
SPLITT Split_263_n653(net36,net120_c1,net202_c1);
SPLITT Split_271_n661(net61,net119_c1,net203_c1);
SPLITT Split_248_n638(net118,net127_c1,net204_c1);
SPLITT Split_256_n646(net113,net125_c1,net205_c1);
SPLITT Split_264_n654(net120,net126_c1,net206_c1);
SPLITT Split_272_n662(net53,net124_c1,net207_c1);
SPLITT Split_280_n670(net78,net123_c1,net208_c1);
SPLITT Split_249_n639(net27,net128_c1,net209_c1);
SPLITT Split_257_n647(net12,net131_c1,net210_c1);
SPLITT Split_265_n655(net52,net130_c1,net211_c1);
SPLITT Split_273_n663(net70,net129_c1,net212_c1);
SPLITT Split_281_n671(net208,net132_c1,net213_c1);
DFFT DFFT_191__FPB_n581(net739,net343,net350_c1);
DFFT DFFT_183__FPB_n573(net393,net344,net348_c1);
DFFT DFFT_175__FPB_n565(net733,net345,net351_c1);
DFFT DFFT_167__FPB_n557(net499,net346,net349_c1);
DFFT DFFT_159__FPB_n549(net392,net347,net352_c1);
SPLITT Split_258_n648(net37,net136_c1,net214_c1);
SPLITT Split_266_n656(net56,net134_c1,net215_c1);
SPLITT Split_274_n664(net84,net133_c1,net216_c1);
SPLITT Split_282_n672(net123,net135_c1,net217_c1);
SPLITT Split_290_n680(net245,net137_c1,net218_c1);
SPLITT Split_259_n649(net11,net141_c1,net219_c1);
SPLITT Split_267_n657(net59,net140_c1,net220_c1);
SPLITT Split_275_n665(net133,net139_c1,net221_c1);
SPLITT Split_283_n673(net82,net138_c1,net222_c1);
SPLITT Split_291_n681(net165,net142_c1,net223_c1);
SPLITT Split_268_n658(net45,net146_c1,net224_c1);
SPLITT Split_276_n666(net88,net145_c1,net225_c1);
SPLITT Split_284_n674(net222,net147_c1,net226_c1);
SPLITT Split_292_n682(net266,net143_c1,net227_c1);
SPLITT Split_269_n659(net54,net151_c1,net229_c1);
SPLITT Split_277_n667(net75,net148_c1,net230_c1);
SPLITT Split_285_n675(net138,net149_c1,net231_c1);
SPLITT Split_293_n683(net227,net152_c1,net232_c1);
SPLITT Split_278_n668(net230,net156_c1,net234_c1);
SPLITT Split_286_n676(net85,net154_c1,net235_c1);
SPLITT Split_294_n684(net143,net155_c1,net236_c1);
SPLITT Split_279_n669(net148,net158_c1,net238_c1);
SPLITT Split_287_n677(net235,net159_c1,net239_c1);
SPLITT Split_295_n685(net267,net157_c1,net240_c1);
SPLITT Split_288_n678(net154,net163_c1,net242_c1);
SPLITT Split_296_n686(net240,net162_c1,net243_c1);
SPLITT Split_289_n679(net81,net165_c1,net245_c1);
SPLITT Split_297_n687(net157,net166_c1,net246_c1);
SPLITT Split_298_n688(net260,net167_c1,net248_c1);
SPLITT Split_299_n689(net167,net170_c1,net250_c1);
DFFT DFFT_192__FPB_n582(net833,net114,net355_c1);
DFFT DFFT_184__FPB_n574(net670,net348,net356_c1);
DFFT DFFT_176__FPB_n566(net823,net200,net357_c1);
DFFT DFFT_168__FPB_n558(net391,net349,net353_c1);
DFFT DFFT_193__FPB_n583(net745,net89,net361_c1);
DFFT DFFT_185__FPB_n575(net390,net246,net358_c1);
DFFT DFFT_177__FPB_n567(net685,net103,net362_c1);
DFFT DFFT_169__FPB_n559(net493,net353,net359_c1);
DFFT DFFT_194__FPB_n584(net723,net87,net365_c1);
DFFT DFFT_186__FPB_n576(net710,net358,net363_c1);
DFFT DFFT_178__FPB_n568(net751,net65,net366_c1);
DFFT DFFT_195__FPB_n585(net706,net98,net368_c1);
DFFT DFFT_187__FPB_n577(net713,net363,net370_c1);
DFFT DFFT_179__FPB_n569(net665,net181,net369_c1);
DFFT DFFT_223_state_obs2(net641,net292,net384_c1);
DFFT DFFT_196__FPB_n586(net707,net368,net372_c1);
DFFT DFFT_188__FPB_n578(net671,net166,net373_c1);
NOTT NOTT_95_n122(net449,net175,net82_c1);
NOTT NOTT_97_n130(net793,net865,net81_c1);
DFFT DFFT_197__FPB_n587(net389,net372,net375_c1);
DFFT DFFT_189__FPB_n579(net711,net373,net376_c1);
DFFT DFFT_216_state_obs1(net627,net299,net383_c1);
DFFT DFFT_98__FPB_n134(net388,net93,net266_c1);
DFFT DFFT_198__FPB_n588(net719,net375,net378_c1);
SPLITT SplitCLK_4_223(net856,net860_c1,net861_c1);
SPLITT SplitCLK_4_224(net857,net858_c1,net859_c1);
SPLITT SplitCLK_6_225(net850,net856_c1,net857_c1);
SPLITT SplitCLK_4_226(net853,net854_c1,net855_c1);
SPLITT SplitCLK_2_227(net851,net852_c1,net853_c1);
SPLITT SplitCLK_0_228(net836,net850_c1,net851_c1);
SPLITT SplitCLK_4_229(net844,net849_c1,net848_c1);
SPLITT SplitCLK_4_230(net845,net847_c1,net846_c1);
SPLITT SplitCLK_6_231(net838,net844_c1,net845_c1);
SPLITT SplitCLK_4_232(net841,net843_c1,net842_c1);
SPLITT SplitCLK_4_233(net839,net840_c1,net841_c1);
SPLITT SplitCLK_6_234(net837,net838_c1,net839_c1);
SPLITT SplitCLK_6_235(net808,net836_c1,net837_c1);
SPLITT SplitCLK_4_236(net830,net835_c1,net834_c1);
SPLITT SplitCLK_4_237(net831,net833_c1,net832_c1);
SPLITT SplitCLK_6_238(net824,net830_c1,net831_c1);
SPLITT SplitCLK_4_239(net827,net828_c1,net829_c1);
SPLITT SplitCLK_4_240(net825,net826_c1,net827_c1);
SPLITT SplitCLK_4_241(net810,net825_c1,net824_c1);
SPLITT SplitCLK_0_242(net818,net823_c1,net822_c1);
SPLITT SplitCLK_4_243(net819,net820_c1,net821_c1);
SPLITT SplitCLK_6_244(net812,net818_c1,net819_c1);
SPLITT SplitCLK_4_245(net815,net817_c1,net816_c1);
SPLITT SplitCLK_2_246(net813,net814_c1,net815_c1);
SPLITT SplitCLK_2_247(net811,net813_c1,net812_c1);
SPLITT SplitCLK_4_248(net809,net811_c1,net810_c1);
SPLITT SplitCLK_0_249(net752,net808_c1,net809_c1);
SPLITT SplitCLK_4_250(net802,net807_c1,net806_c1);
SPLITT SplitCLK_4_251(net803,net804_c1,net805_c1);
SPLITT SplitCLK_6_252(net796,net802_c1,net803_c1);
SPLITT SplitCLK_4_253(net799,net800_c1,net801_c1);
SPLITT SplitCLK_0_254(net797,net798_c1,net799_c1);
SPLITT SplitCLK_6_255(net782,net797_c1,net796_c1);
SPLITT SplitCLK_4_256(net790,net794_c1,net795_c1);
SPLITT SplitCLK_4_257(net791,net792_c1,net793_c1);
SPLITT SplitCLK_6_258(net784,net790_c1,net791_c1);
SPLITT SplitCLK_4_259(net787,net788_c1,net789_c1);
SPLITT SplitCLK_4_260(net785,net786_c1,net787_c1);
SPLITT SplitCLK_6_261(net783,net785_c1,net784_c1);
SPLITT SplitCLK_6_262(net754,net782_c1,net783_c1);
SPLITT SplitCLK_4_263(net776,net781_c1,net780_c1);
SPLITT SplitCLK_4_264(net777,net779_c1,net778_c1);
SPLITT SplitCLK_6_265(net770,net776_c1,net777_c1);
SPLITT SplitCLK_4_266(net773,net775_c1,net774_c1);
SPLITT SplitCLK_4_267(net771,net772_c1,net773_c1);
SPLITT SplitCLK_0_268(net756,net770_c1,net771_c1);
SPLITT SplitCLK_4_269(net764,net769_c1,net768_c1);
SPLITT SplitCLK_4_270(net765,net767_c1,net766_c1);
SPLITT SplitCLK_6_271(net758,net764_c1,net765_c1);
SPLITT SplitCLK_4_272(net761,net762_c1,net763_c1);
SPLITT SplitCLK_4_273(net759,net760_c1,net761_c1);
SPLITT SplitCLK_2_274(net757,net759_c1,net758_c1);
SPLITT SplitCLK_4_275(net755,net757_c1,net756_c1);
SPLITT SplitCLK_2_276(net753,net755_c1,net754_c1);
SPLITT SplitCLK_6_277(net642,net752_c1,net753_c1);
SPLITT SplitCLK_4_278(net746,net751_c1,net750_c1);
SPLITT SplitCLK_4_279(net747,net748_c1,net749_c1);
SPLITT SplitCLK_4_280(net740,net747_c1,net746_c1);
SPLITT SplitCLK_4_281(net743,net745_c1,net744_c1);
SPLITT SplitCLK_2_282(net741,net743_c1,net742_c1);
SPLITT SplitCLK_4_283(net726,net741_c1,net740_c1);
SPLITT SplitCLK_4_284(net734,net739_c1,net738_c1);
SPLITT SplitCLK_4_285(net735,net736_c1,net737_c1);
SPLITT SplitCLK_6_286(net728,net734_c1,net735_c1);
SPLITT SplitCLK_4_287(net731,net733_c1,net732_c1);
SPLITT SplitCLK_4_288(net729,net730_c1,net731_c1);
SPLITT SplitCLK_2_289(net727,net729_c1,net728_c1);
SPLITT SplitCLK_6_290(net698,net726_c1,net727_c1);
SPLITT SplitCLK_4_291(net720,net724_c1,net725_c1);
SPLITT SplitCLK_4_292(net721,net723_c1,net722_c1);
SPLITT SplitCLK_4_293(net714,net721_c1,net720_c1);
SPLITT SplitCLK_4_294(net717,net718_c1,net719_c1);
SPLITT SplitCLK_4_295(net715,net716_c1,net717_c1);
SPLITT SplitCLK_0_296(net700,net714_c1,net715_c1);
SPLITT SplitCLK_4_297(net708,net712_c1,net713_c1);
SPLITT SplitCLK_4_298(net709,net711_c1,net710_c1);
SPLITT SplitCLK_4_299(net702,net709_c1,net708_c1);
SPLITT SplitCLK_4_300(net705,net706_c1,net707_c1);
SPLITT SplitCLK_4_301(net703,net704_c1,net705_c1);
SPLITT SplitCLK_2_302(net701,net702_c1,net703_c1);
SPLITT SplitCLK_4_303(net699,net701_c1,net700_c1);
SPLITT SplitCLK_0_304(net644,net698_c1,net699_c1);
SPLITT SplitCLK_4_305(net692,net696_c1,net697_c1);
SPLITT SplitCLK_0_306(net693,net694_c1,net695_c1);
SPLITT SplitCLK_0_307(net686,net693_c1,net692_c1);
SPLITT SplitCLK_4_308(net689,net691_c1,net690_c1);
SPLITT SplitCLK_2_309(net687,net689_c1,net688_c1);
SPLITT SplitCLK_4_310(net672,net687_c1,net686_c1);
SPLITT SplitCLK_4_311(net680,net684_c1,net685_c1);
SPLITT SplitCLK_0_312(net681,net682_c1,net683_c1);
SPLITT SplitCLK_6_313(net674,net680_c1,net681_c1);
SPLITT SplitCLK_4_314(net677,net678_c1,net679_c1);
SPLITT SplitCLK_4_315(net675,net676_c1,net677_c1);
SPLITT SplitCLK_2_316(net673,net674_c1,net675_c1);
SPLITT SplitCLK_6_317(net646,net672_c1,net673_c1);
SPLITT SplitCLK_4_318(net666,net670_c1,net671_c1);
SPLITT SplitCLK_4_319(net667,net669_c1,net668_c1);
SPLITT SplitCLK_6_320(net660,net666_c1,net667_c1);
SPLITT SplitCLK_4_321(net663,net665_c1,net664_c1);
SPLITT SplitCLK_4_322(net661,net662_c1,net663_c1);
SPLITT SplitCLK_0_323(net648,net660_c1,net661_c1);
SPLITT SplitCLK_4_324(net657,net659_c1,net658_c1);
SPLITT SplitCLK_2_325(net650,net657_c1,net656_c1);
SPLITT SplitCLK_4_326(net653,net655_c1,net654_c1);
SPLITT SplitCLK_4_327(net651,net652_c1,net653_c1);
SPLITT SplitCLK_6_328(net649,net651_c1,net650_c1);
SPLITT SplitCLK_4_329(net647,net649_c1,net648_c1);
SPLITT SplitCLK_2_330(net645,net647_c1,net646_c1);
SPLITT SplitCLK_4_331(net643,net645_c1,net644_c1);
SPLITT SplitCLK_0_332(net386,net642_c1,net643_c1);
SPLITT SplitCLK_4_333(net636,net641_c1,net640_c1);
SPLITT SplitCLK_0_334(net637,net638_c1,net639_c1);
SPLITT SplitCLK_0_335(net630,net637_c1,net636_c1);
SPLITT SplitCLK_4_336(net633,net634_c1,net635_c1);
SPLITT SplitCLK_6_337(net631,net633_c1,net632_c1);
SPLITT SplitCLK_4_338(net616,net631_c1,net630_c1);
SPLITT SplitCLK_4_339(net624,net629_c1,net628_c1);
SPLITT SplitCLK_0_340(net625,net626_c1,net627_c1);
SPLITT SplitCLK_0_341(net618,net625_c1,net624_c1);
SPLITT SplitCLK_4_342(net621,net622_c1,net623_c1);
SPLITT SplitCLK_2_343(net619,net620_c1,net621_c1);
SPLITT SplitCLK_2_344(net617,net618_c1,net619_c1);
SPLITT SplitCLK_6_345(net588,net616_c1,net617_c1);
SPLITT SplitCLK_4_346(net610,net614_c1,net615_c1);
SPLITT SplitCLK_0_347(net611,net612_c1,net613_c1);
SPLITT SplitCLK_0_348(net604,net611_c1,net610_c1);
SPLITT SplitCLK_4_349(net607,net609_c1,net608_c1);
SPLITT SplitCLK_2_350(net605,net606_c1,net607_c1);
SPLITT SplitCLK_4_351(net590,net605_c1,net604_c1);
SPLITT SplitCLK_4_352(net598,net603_c1,net602_c1);
SPLITT SplitCLK_0_353(net599,net601_c1,net600_c1);
SPLITT SplitCLK_6_354(net592,net598_c1,net599_c1);
SPLITT SplitCLK_4_355(net595,net597_c1,net596_c1);
SPLITT SplitCLK_4_356(net593,net594_c1,net595_c1);
SPLITT SplitCLK_2_357(net591,net593_c1,net592_c1);
SPLITT SplitCLK_4_358(net589,net591_c1,net590_c1);
SPLITT SplitCLK_6_359(net532,net589_c1,net588_c1);
SPLITT SplitCLK_4_360(net582,net587_c1,net586_c1);
SPLITT SplitCLK_0_361(net583,net584_c1,net585_c1);
SPLITT SplitCLK_0_362(net576,net583_c1,net582_c1);
SPLITT SplitCLK_4_363(net579,net581_c1,net580_c1);
SPLITT SplitCLK_0_364(net577,net578_c1,net579_c1);
SPLITT SplitCLK_4_365(net562,net576_c1,net577_c1);
SPLITT SplitCLK_4_366(net570,net575_c1,net574_c1);
SPLITT SplitCLK_4_367(net571,net572_c1,net573_c1);
SPLITT SplitCLK_4_368(net564,net571_c1,net570_c1);
SPLITT SplitCLK_4_369(net567,net569_c1,net568_c1);
SPLITT SplitCLK_2_370(net565,net566_c1,net567_c1);
SPLITT SplitCLK_2_371(net563,net565_c1,net564_c1);
SPLITT SplitCLK_6_372(net534,net562_c1,net563_c1);
SPLITT SplitCLK_4_373(net556,net561_c1,net560_c1);
SPLITT SplitCLK_0_374(net557,net559_c1,net558_c1);
SPLITT SplitCLK_0_375(net550,net557_c1,net556_c1);
SPLITT SplitCLK_4_376(net553,net554_c1,net555_c1);
SPLITT SplitCLK_4_377(net551,net552_c1,net553_c1);
SPLITT SplitCLK_4_378(net536,net550_c1,net551_c1);
SPLITT SplitCLK_4_379(net544,net549_c1,net548_c1);
SPLITT SplitCLK_4_380(net545,net546_c1,net547_c1);
SPLITT SplitCLK_6_381(net538,net544_c1,net545_c1);
SPLITT SplitCLK_4_382(net541,net543_c1,net542_c1);
SPLITT SplitCLK_4_383(net539,net540_c1,net541_c1);
SPLITT SplitCLK_2_384(net537,net539_c1,net538_c1);
SPLITT SplitCLK_4_385(net535,net537_c1,net536_c1);
SPLITT SplitCLK_2_386(net533,net535_c1,net534_c1);
SPLITT SplitCLK_6_387(net422,net532_c1,net533_c1);
SPLITT SplitCLK_4_388(net526,net531_c1,net530_c1);
SPLITT SplitCLK_4_389(net527,net528_c1,net529_c1);
SPLITT SplitCLK_6_390(net520,net526_c1,net527_c1);
SPLITT SplitCLK_4_391(net523,net524_c1,net525_c1);
SPLITT SplitCLK_4_392(net521,net522_c1,net523_c1);
SPLITT SplitCLK_0_393(net506,net520_c1,net521_c1);
SPLITT SplitCLK_4_394(net514,net518_c1,net519_c1);
SPLITT SplitCLK_4_395(net515,net517_c1,net516_c1);
SPLITT SplitCLK_2_396(net508,net514_c1,net515_c1);
SPLITT SplitCLK_4_397(net511,net513_c1,net512_c1);
SPLITT SplitCLK_2_398(net509,net510_c1,net511_c1);
SPLITT SplitCLK_2_399(net507,net509_c1,net508_c1);
SPLITT SplitCLK_6_400(net478,net506_c1,net507_c1);
SPLITT SplitCLK_4_401(net500,net504_c1,net505_c1);
SPLITT SplitCLK_4_402(net501,net503_c1,net502_c1);
SPLITT SplitCLK_6_403(net494,net500_c1,net501_c1);
SPLITT SplitCLK_4_404(net497,net499_c1,net498_c1);
SPLITT SplitCLK_4_405(net495,net496_c1,net497_c1);
SPLITT SplitCLK_4_406(net480,net494_c1,net495_c1);
SPLITT SplitCLK_0_407(net488,net492_c1,net493_c1);
SPLITT SplitCLK_4_408(net489,net490_c1,net491_c1);
SPLITT SplitCLK_4_409(net482,net489_c1,net488_c1);
SPLITT SplitCLK_4_410(net485,net486_c1,net487_c1);
SPLITT SplitCLK_2_411(net483,net485_c1,net484_c1);
SPLITT SplitCLK_6_412(net481,net482_c1,net483_c1);
SPLITT SplitCLK_4_413(net479,net481_c1,net480_c1);
SPLITT SplitCLK_0_414(net424,net478_c1,net479_c1);
SPLITT SplitCLK_4_415(net472,net477_c1,net476_c1);
SPLITT SplitCLK_4_416(net473,net475_c1,net474_c1);
SPLITT SplitCLK_4_417(net466,net473_c1,net472_c1);
SPLITT SplitCLK_4_418(net469,net470_c1,net471_c1);
SPLITT SplitCLK_4_419(net467,net468_c1,net469_c1);
SPLITT SplitCLK_0_420(net452,net466_c1,net467_c1);
SPLITT SplitCLK_4_421(net460,net464_c1,net465_c1);
SPLITT SplitCLK_4_422(net461,net462_c1,net463_c1);
SPLITT SplitCLK_2_423(net454,net460_c1,net461_c1);
SPLITT SplitCLK_4_424(net457,net459_c1,net458_c1);
SPLITT SplitCLK_4_425(net455,net456_c1,net457_c1);
SPLITT SplitCLK_2_426(net453,net455_c1,net454_c1);
SPLITT SplitCLK_6_427(net426,net452_c1,net453_c1);
SPLITT SplitCLK_4_428(net446,net450_c1,net451_c1);
SPLITT SplitCLK_4_429(net447,net449_c1,net448_c1);
SPLITT SplitCLK_0_430(net440,net446_c1,net447_c1);
SPLITT SplitCLK_4_431(net443,net445_c1,net444_c1);
SPLITT SplitCLK_4_432(net441,net442_c1,net443_c1);
SPLITT SplitCLK_0_433(net428,net440_c1,net441_c1);
SPLITT SplitCLK_4_434(net437,net439_c1,net438_c1);
SPLITT SplitCLK_2_435(net430,net437_c1,net436_c1);
SPLITT SplitCLK_4_436(net433,net435_c1,net434_c1);
SPLITT SplitCLK_2_437(net431,net432_c1,net433_c1);
SPLITT SplitCLK_2_438(net429,net431_c1,net430_c1);
SPLITT SplitCLK_4_439(net427,net429_c1,net428_c1);
SPLITT SplitCLK_2_440(net425,net427_c1,net426_c1);
SPLITT SplitCLK_4_441(net423,net425_c1,net424_c1);
SPLITT SplitCLK_2_442(net387,net423_c1,net422_c1);
wire dummy0;
SPLITT SplitCLK_2_443(net578,net421_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_2_444(net772,net420_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_445(net594,net419_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_4_446(net552,net418_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_447(net456,net417_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_2_448(net522,net416_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_2_449(net826,net415_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_2_450(net760,net414_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_2_451(net676,net413_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_2_452(net814,net412_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_2_453(net620,net411_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_2_454(net798,net410_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_2_455(net786,net409_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_2_456(net742,net408_c1,dummy13);
wire dummy14;
SPLITT SplitCLK_2_457(net688,net407_c1,dummy14);
wire dummy15;
SPLITT SplitCLK_4_458(net632,net406_c1,dummy15);
wire dummy16;
SPLITT SplitCLK_4_459(net540,net405_c1,dummy16);
wire dummy17;
SPLITT SplitCLK_2_460(net852,net404_c1,dummy17);
wire dummy18;
SPLITT SplitCLK_2_461(net436,net403_c1,dummy18);
wire dummy19;
SPLITT SplitCLK_2_462(net566,net402_c1,dummy19);
wire dummy20;
SPLITT SplitCLK_2_463(net606,net401_c1,dummy20);
wire dummy21;
SPLITT SplitCLK_2_464(net468,net400_c1,dummy21);
wire dummy22;
SPLITT SplitCLK_2_465(net510,net399_c1,dummy22);
wire dummy23;
SPLITT SplitCLK_2_466(net656,net398_c1,dummy23);
wire dummy24;
SPLITT SplitCLK_2_467(net840,net397_c1,dummy24);
wire dummy25;
SPLITT SplitCLK_2_468(net442,net396_c1,dummy25);
wire dummy26;
SPLITT SplitCLK_2_469(net432,net395_c1,dummy26);
wire dummy27;
SPLITT SplitCLK_2_470(net730,net394_c1,dummy27);
wire dummy28;
SPLITT SplitCLK_2_471(net662,net393_c1,dummy28);
wire dummy29;
SPLITT SplitCLK_2_472(net652,net392_c1,dummy29);
wire dummy30;
SPLITT SplitCLK_2_473(net496,net391_c1,dummy30);
wire dummy31;
SPLITT SplitCLK_2_474(net704,net390_c1,dummy31);
wire dummy32;
SPLITT SplitCLK_2_475(net716,net389_c1,dummy32);
wire dummy33;
SPLITT SplitCLK_2_476(net484,net388_c1,dummy33);
SPLITT SplitCLK_0_477(net862,net386_c1,net387_c1);
wire dummy34;
SPLITT Split_HOLD_566(net308,dummy34,net863_c1);
wire dummy35;
SPLITT Split_HOLD_567(net287,dummy35,net864_c1);
wire dummy36;
SPLITT Split_HOLD_568(net265,dummy36,net865_c1);
wire dummy37;
SPLITT Split_HOLD_569(net283,dummy37,net866_c1);
wire dummy38;
SPLITT Split_HOLD_570(net367,dummy38,net867_c1);
wire dummy39;
SPLITT Split_HOLD_571(net273,dummy39,net868_c1);
INTERCONNECT TMS_Pad_Split_230_n620(TMS_Pad,net0);
INTERCONNECT OR2T_16_n40_DFFT_103__PIPL_n139(net1_c1,net1);
INTERCONNECT NOTT_8_n32_Split_232_n622(net2_c1,net2);
INTERCONNECT NOTT_17_n41_Split_240_n630(net3_c1,net3);
INTERCONNECT NOTT_9_n33_DFFT_100__PIPL_n136(net4_c1,net4);
INTERCONNECT AND2T_26_n50_OR2T_27_n51(net5_c1,net5);
INTERCONNECT NOTT_18_n42_Split_243_n633(net6_c1,net6);
INTERCONNECT NOTT_10_n34_Split_235_n625(net7_c1,net7);
INTERCONNECT OR2T_27_n51_OR2T_28_n52(net8_c1,net8);
INTERCONNECT AND2T_19_n43_Split_244_n634(net9_c1,net9);
INTERCONNECT NOTT_11_n35_DFFT_101__PIPL_n137(net10_c1,net10);
INTERCONNECT AND2T_36_n60_Split_259_n649(net11_c1,net11);
INTERCONNECT OR2T_28_n52_Split_257_n647(net12_c1,net12);
INTERCONNECT AND2T_20_n44_DFFT_121__FPB_n511(net13_c1,net13);
INTERCONNECT NOTT_12_n36_AND2T_94_n121(net14_c1,net14);
INTERCONNECT OR2T_37_n61_OR2T_38_n62(net15_c1,net15);
INTERCONNECT AND2T_29_n53_DFFT_143__FPB_n533(net16_c1,net16);
INTERCONNECT AND2T_21_n45_Split_247_n637(net17_c1,net17);
INTERCONNECT NOTT_13_n37_DFFT_102__PIPL_n138(net18_c1,net18);
INTERCONNECT OR2T_46_n70_OR2T_49_n73(net19_c1,net19);
INTERCONNECT OR2T_38_n62_AND2T_39_n63(net20_c1,net20);
INTERCONNECT AND2T_30_n54_AND2T_77_n101(net21_c1,net21);
INTERCONNECT AND2T_22_n46_DFFT_120__FPB_n510(net22_c1,net22);
INTERCONNECT AND2T_14_n38_Split_238_n628(net23_c1,net23);
INTERCONNECT AND2T_47_n71_DFFT_141__FPB_n531(net24_c1,net24);
INTERCONNECT AND2T_39_n63_OR2T_51_n75(net25_c1,net25);
INTERCONNECT AND2T_31_n55_OR2T_33_n57(net26_c1,net26);
INTERCONNECT NOTT_23_n47_Split_249_n639(net27_c1,net27);
INTERCONNECT AND2T_15_n39_Split_239_n629(net28_c1,net28);
INTERCONNECT AND2T_56_n80_OR2T_68_n92(net29_c1,net29);
INTERCONNECT XOR2T_48_n72_AND2T_47_n71(net30_c1,net30);
INTERCONNECT AND2T_40_n64_Split_260_n650(net31_c1,net31);
INTERCONNECT AND2T_32_n56_OR2T_33_n57(net32_c1,net32);
INTERCONNECT AND2T_24_n48_Split_251_n641(net33_c1,net33);
INTERCONNECT AND2T_57_n81_OR2T_59_n83(net34_c1,net34);
INTERCONNECT OR2T_49_n73_OR2T_50_n74(net35_c1,net35);
INTERCONNECT AND2T_41_n65_Split_263_n653(net36_c1,net36);
INTERCONNECT OR2T_33_n57_Split_258_n648(net37_c1,net37);
INTERCONNECT AND2T_25_n49_Split_254_n644(net38_c1,net38);
INTERCONNECT OR2T_66_n90_OR2T_67_n91(net39_c1,net39);
INTERCONNECT AND2T_58_n82_OR2T_59_n83(net40_c1,net40);
INTERCONNECT OR2T_50_n74_OR2T_51_n75(net41_c1,net41);
INTERCONNECT AND2T_42_n66_DFFT_142__FPB_n532(net42_c1,net42);
INTERCONNECT OR2T_34_n58_AND2T_39_n63(net43_c1,net43);
INTERCONNECT OR2T_67_n91_OR2T_68_n92(net44_c1,net44);
INTERCONNECT OR2T_59_n83_Split_268_n658(net45_c1,net45);
INTERCONNECT OR2T_51_n75_OR2T_52_n76(net46_c1,net46);
INTERCONNECT AND2T_43_n67_AND2T_44_n68(net47_c1,net47);
INTERCONNECT AND2T_35_n59_DFFT_134__FPB_n524(net48_c1,net48);
INTERCONNECT OR2T_68_n92_AND2T_69_n93(net49_c1,net49);
INTERCONNECT AND2T_60_n84_DFFT_164__FPB_n554(net50_c1,net50);
INTERCONNECT OR2T_52_n76_AND2T_53_n77(net51_c1,net51);
INTERCONNECT AND2T_44_n68_Split_265_n655(net52_c1,net52);
INTERCONNECT AND2T_69_n93_Split_272_n662(net53_c1,net53);
INTERCONNECT AND2T_61_n85_Split_269_n659(net54_c1,net54);
INTERCONNECT AND2T_53_n77_DFFT_104__FBL_n494(net55_c1,net55);
INTERCONNECT AND2T_45_n69_Split_266_n656(net56_c1,net56);
INTERCONNECT AND2T_70_n94_AND2T_71_n95(net57_c1,net57);
INTERCONNECT AND2T_62_n86_Split_270_n660(net58_c1,net58);
INTERCONNECT OR2T_54_n78_Split_267_n657(net59_c1,net59);
INTERCONNECT AND2T_71_n95_OR2T_72_n96(net60_c1,net60);
INTERCONNECT AND2T_63_n87_Split_271_n661(net61_c1,net61);
INTERCONNECT OR2T_55_n79_AND2T_56_n80(net62_c1,net62);
INTERCONNECT OR2T_72_n96_OR2T_73_n97(net63_c1,net63);
INTERCONNECT OR2T_64_n88_OR2T_65_n89(net64_c1,net64);
INTERCONNECT OR2T_73_n97_DFFT_178__FPB_n568(net65_c1,net65);
INTERCONNECT OR2T_65_n89_OR2T_66_n90(net66_c1,net66);
INTERCONNECT AND2T_74_n98_OR2T_75_n99(net67_c1,net67);
INTERCONNECT OR2T_75_n99_OR2T_80_n104(net68_c1,net68);
INTERCONNECT AND2T_76_n100_OR2T_79_n103(net69_c1,net69);
INTERCONNECT AND2T_77_n101_Split_273_n663(net70_c1,net70);
INTERCONNECT AND2T_86_n110_OR2T_88_n112(net71_c1,net71);
INTERCONNECT AND2T_78_n102_OR2T_79_n103(net72_c1,net72);
INTERCONNECT OR2T_87_n111_AND2T_86_n110(net73_c1,net73);
INTERCONNECT OR2T_79_n103_OR2T_80_n104(net74_c1,net74);
INTERCONNECT AND2T_93_n120_Split_277_n667(net75_c1,net75);
INTERCONNECT OR2T_88_n112_OR2T_89_n113(net76_c1,net76);
INTERCONNECT OR2T_80_n104_OR2T_81_n105(net77_c1,net77);
INTERCONNECT AND2T_94_n121_Split_280_n670(net78_c1,net78);
INTERCONNECT OR2T_89_n113_OR2T_90_n114(net79_c1,net79);
INTERCONNECT OR2T_81_n105_AND2T_82_n106(net80_c1,net80);
INTERCONNECT NOTT_97_n130_Split_289_n679(net81_c1,net81);
INTERCONNECT NOTT_95_n122_Split_283_n673(net82_c1,net82);
INTERCONNECT OR2T_90_n114_OR2T_91_n115(net83_c1,net83);
INTERCONNECT AND2T_82_n106_Split_274_n664(net84_c1,net84);
INTERCONNECT AND2T_96_n123_Split_286_n676(net85_c1,net85);
INTERCONNECT OR2T_91_n115_AND2T_92_n116(net86_c1,net86);
INTERCONNECT AND2T_83_n107_DFFT_194__FPB_n584(net87_c1,net87);
INTERCONNECT AND2T_92_n116_Split_276_n666(net88_c1,net88);
INTERCONNECT AND2T_84_n108_DFFT_193__FPB_n583(net89_c1,net89);
INTERCONNECT AND2T_85_n109_OR2T_88_n112(net90_c1,net90);
INTERCONNECT Split_230_n620_Split_231_n621(net91_c1,net91);
INTERCONNECT Split_310_n700_DFFT_126__FPB_n516(net92_c1,net92);
INTERCONNECT Split_231_n621_DFFT_98__FPB_n134(net93_c1,net93);
INTERCONNECT Split_240_n630_Split_242_n632(net94_c1,net94);
INTERCONNECT Split_232_n622_Split_234_n624(net95_c1,net95);
INTERCONNECT Split_241_n631_DFFT_165__FPB_n555(net96_c1,net96);
INTERCONNECT Split_233_n623_AND2T_19_n43(net97_c1,net97);
INTERCONNECT Split_242_n632_DFFT_195__FPB_n585(net98_c1,net98);
INTERCONNECT Split_234_n624_OR2T_87_n111(net99_c1,net99);
INTERCONNECT Split_250_n640_AND2T_30_n54(net100_c1,net100);
INTERCONNECT Split_251_n641_Split_253_n643(net101_c1,net101);
INTERCONNECT Split_235_n625_Split_237_n627(net102_c1,net102);
INTERCONNECT Split_243_n633_DFFT_177__FPB_n567(net103_c1,net103);
INTERCONNECT Split_260_n650_Split_262_n652(net104_c1,net104);
INTERCONNECT Split_244_n634_Split_246_n636(net105_c1,net105);
INTERCONNECT Split_252_n642_AND2T_32_n56(net106_c1,net106);
INTERCONNECT Split_236_n626_AND2T_19_n43(net107_c1,net107);
INTERCONNECT TRST_Pad_NOTT_17_n41(TRST_Pad,net108);
INTERCONNECT Split_261_n651_AND2T_47_n71(net109_c1,net109);
INTERCONNECT Split_253_n643_AND2T_57_n81(net110_c1,net110);
INTERCONNECT Split_237_n627_OR2T_87_n111(net111_c1,net111);
INTERCONNECT Split_245_n635_AND2T_31_n55(net112_c1,net112);
INTERCONNECT Split_254_n644_Split_256_n646(net113_c1,net113);
INTERCONNECT Split_238_n628_DFFT_192__FPB_n582(net114_c1,net114);
INTERCONNECT Split_270_n660_DFFT_163__FPB_n553(net115_c1,net115);
INTERCONNECT Split_262_n652_AND2T_63_n87(net116_c1,net116);
INTERCONNECT Split_246_n636_AND2T_45_n69(net117_c1,net117);
INTERCONNECT Split_247_n637_Split_248_n638(net118_c1,net118);
INTERCONNECT Split_271_n661_DFFT_162__FPB_n552(net119_c1,net119);
INTERCONNECT Split_263_n653_Split_264_n654(net120_c1,net120);
INTERCONNECT Split_239_n629_AND2T_85_n109(net121_c1,net121);
INTERCONNECT Split_255_n645_AND2T_36_n60(net122_c1,net122);
INTERCONNECT Split_280_n670_Split_282_n672(net123_c1,net123);
INTERCONNECT Split_272_n662_DFFT_108__FBL_n498(net124_c1,net124);
INTERCONNECT Split_256_n646_AND2T_61_n85(net125_c1,net125);
INTERCONNECT Split_264_n654_OR2T_64_n88(net126_c1,net126);
INTERCONNECT Split_248_n638_DFFT_127__FPB_n517(net127_c1,net127);
INTERCONNECT Split_249_n639_Split_250_n640(net128_c1,net128);
INTERCONNECT Split_273_n663_AND2T_84_n108(net129_c1,net129);
INTERCONNECT Split_265_n655_OR2T_64_n88(net130_c1,net130);
INTERCONNECT Split_257_n647_OR2T_55_n79(net131_c1,net131);
INTERCONNECT Split_281_n671_AND2T_20_n44(net132_c1,net132);
INTERCONNECT Split_274_n664_Split_275_n665(net133_c1,net133);
INTERCONNECT Split_266_n656_OR2T_54_n78(net134_c1,net134);
INTERCONNECT Split_282_n672_DFFT_160__FPB_n550(net135_c1,net135);
INTERCONNECT Split_258_n648_OR2T_73_n97(net136_c1,net136);
INTERCONNECT Split_290_n680_AND2T_15_n39(net137_c1,net137);
INTERCONNECT Split_283_n673_Split_285_n675(net138_c1,net138);
INTERCONNECT Split_275_n665_DFFT_114__FPB_n504(net139_c1,net139);
INTERCONNECT Split_267_n657_DFFT_151__FPB_n541(net140_c1,net140);
INTERCONNECT Split_259_n649_OR2T_54_n78(net141_c1,net141);
INTERCONNECT Split_291_n681_XOR2T_48_n72(net142_c1,net142);
INTERCONNECT Split_292_n682_Split_294_n684(net143_c1,net143);
INTERCONNECT Split_300_n690_DFFT_190__FPB_n580(net144_c1,net144);
INTERCONNECT Split_276_n666_DFFT_115__FPB_n505(net145_c1,net145);
INTERCONNECT Split_268_n658_AND2T_83_n107(net146_c1,net146);
INTERCONNECT Split_284_n674_DFFT_122__FPB_n512(net147_c1,net147);
INTERCONNECT Split_277_n667_Split_279_n669(net148_c1,net148);
INTERCONNECT Split_285_n675_DFFT_157__FPB_n547(net149_c1,net149);
INTERCONNECT Split_301_n691_DFFT_201__FPB_n591(net150_c1,net150);
INTERCONNECT Split_269_n659_AND2T_74_n98(net151_c1,net151);
INTERCONNECT Split_293_n683_DFFT_132__FPB_n522(net152_c1,net152);
INTERCONNECT Split_302_n692_Split_304_n694(net153_c1,net153);
INTERCONNECT Split_286_n676_Split_288_n678(net154_c1,net154);
INTERCONNECT Split_294_n684_DFFT_152__FPB_n542(net155_c1,net155);
INTERCONNECT Split_278_n668_DFFT_118__FPB_n508(net156_c1,net156);
INTERCONNECT Split_295_n685_Split_297_n687(net157_c1,net157);
INTERCONNECT Split_279_n669_DFFT_139__FPB_n529(net158_c1,net158);
INTERCONNECT Split_287_n677_AND2T_41_n65(net159_c1,net159);
INTERCONNECT Split_303_n693_AND2T_21_n45(net160_c1,net160);
INTERCONNECT Split_304_n694_DFFT_138__FPB_n528(net161_c1,net161);
INTERCONNECT Split_296_n686_DFFT_174__FPB_n564(net162_c1,net162);
INTERCONNECT Split_288_n678_DFFT_173__FPB_n563(net163_c1,net163);
INTERCONNECT Split_305_n695_Split_307_n697(net164_c1,net164);
INTERCONNECT Split_289_n679_Split_291_n681(net165_c1,net165);
INTERCONNECT Split_297_n687_DFFT_188__FPB_n578(net166_c1,net166);
INTERCONNECT Split_298_n688_Split_299_n689(net167_c1,net167);
INTERCONNECT Split_306_n696_NOTT_23_n47(net168_c1,net168);
INTERCONNECT Split_307_n697_DFFT_140__FPB_n530(net169_c1,net169);
INTERCONNECT Split_299_n689_AND2T_21_n45(net170_c1,net170);
INTERCONNECT Split_308_n698_Split_310_n700(net171_c1,net171);
INTERCONNECT Split_309_n699_AND2T_14_n38(net172_c1,net172);
INTERCONNECT Split_230_n620_DFFT_99__FPB_n135(net173_c1,net173);
INTERCONNECT Split_310_n700_AND2T_93_n120(net174_c1,net174);
INTERCONNECT Split_231_n621_NOTT_95_n122(net175_c1,net175);
INTERCONNECT Split_232_n622_Split_233_n623(net176_c1,net176);
INTERCONNECT Split_240_n630_Split_241_n631(net177_c1,net177);
INTERCONNECT Split_233_n623_NOTT_9_n33(net178_c1,net178);
INTERCONNECT Split_241_n631_DFFT_144__FPB_n534(net179_c1,net179);
INTERCONNECT Split_234_n624_AND2T_40_n64(net180_c1,net180);
INTERCONNECT Split_242_n632_DFFT_179__FPB_n569(net181_c1,net181);
INTERCONNECT Split_250_n640_AND2T_24_n48(net182_c1,net182);
INTERCONNECT Split_235_n625_Split_236_n626(net183_c1,net183);
INTERCONNECT Split_243_n633_AND2T_61_n85(net184_c1,net184);
INTERCONNECT Split_251_n641_Split_252_n642(net185_c1,net185);
INTERCONNECT Split_236_n626_NOTT_11_n35(net186_c1,net186);
INTERCONNECT Split_244_n634_Split_245_n635(net187_c1,net187);
INTERCONNECT Split_252_n642_AND2T_26_n50(net188_c1,net188);
INTERCONNECT Split_260_n650_Split_261_n651(net189_c1,net189);
INTERCONNECT Split_237_n627_AND2T_25_n49(net190_c1,net190);
INTERCONNECT Split_245_n635_AND2T_20_n44(net191_c1,net191);
INTERCONNECT Split_253_n643_AND2T_35_n59(net192_c1,net192);
INTERCONNECT Split_261_n651_AND2T_41_n65(net193_c1,net193);
INTERCONNECT Split_238_n628_DFFT_161__FPB_n551(net194_c1,net194);
INTERCONNECT Split_246_n636_AND2T_35_n59(net195_c1,net195);
INTERCONNECT Split_254_n644_Split_255_n645(net196_c1,net196);
INTERCONNECT Split_262_n652_AND2T_57_n81(net197_c1,net197);
INTERCONNECT Split_270_n660_OR2T_89_n113(net198_c1,net198);
INTERCONNECT Split_239_n629_AND2T_71_n95(net199_c1,net199);
INTERCONNECT Split_247_n637_DFFT_176__FPB_n566(net200_c1,net200);
INTERCONNECT Split_255_n645_AND2T_26_n50(net201_c1,net201);
INTERCONNECT Split_263_n653_OR2T_72_n96(net202_c1,net202);
INTERCONNECT Split_271_n661_AND2T_76_n100(net203_c1,net203);
INTERCONNECT Split_248_n638_AND2T_22_n46(net204_c1,net204);
INTERCONNECT Split_256_n646_AND2T_58_n82(net205_c1,net205);
INTERCONNECT Split_264_n654_AND2T_42_n66(net206_c1,net206);
INTERCONNECT Split_272_n662_DFFT_105__FBL_n495(net207_c1,net207);
INTERCONNECT Split_280_n670_Split_281_n671(net208_c1,net208);
INTERCONNECT Split_249_n639_AND2T_96_n123(net209_c1,net209);
INTERCONNECT Split_257_n647_AND2T_29_n53(net210_c1,net210);
INTERCONNECT Split_265_n655_OR2T_46_n70(net211_c1,net211);
INTERCONNECT Split_273_n663_AND2T_78_n102(net212_c1,net212);
INTERCONNECT Split_281_n671_OR2T_16_n40(net213_c1,net213);
INTERCONNECT Split_258_n648_OR2T_34_n58(net214_c1,net214);
INTERCONNECT Split_266_n656_OR2T_46_n70(net215_c1,net215);
INTERCONNECT Split_274_n664_DFFT_116__FPB_n506(net216_c1,net216);
INTERCONNECT Split_282_n672_AND2T_44_n68(net217_c1,net217);
INTERCONNECT Split_290_n680_NOTT_13_n37(net218_c1,net218);
INTERCONNECT Split_259_n649_OR2T_37_n61(net219_c1,net219);
INTERCONNECT Split_267_n657_OR2T_75_n99(net220_c1,net220);
INTERCONNECT Split_275_n665_DFFT_112__FPB_n502(net221_c1,net221);
INTERCONNECT Split_283_n673_Split_284_n674(net222_c1,net222);
INTERCONNECT Split_291_n681_AND2T_24_n48(net223_c1,net223);
INTERCONNECT Split_268_n658_AND2T_60_n84(net224_c1,net224);
INTERCONNECT Split_276_n666_DFFT_113__FPB_n503(net225_c1,net225);
INTERCONNECT Split_284_n674_AND2T_43_n67(net226_c1,net226);
INTERCONNECT Split_292_n682_Split_293_n683(net227_c1,net227);
INTERCONNECT Split_300_n690_DFFT_172__FPB_n562(net228_c1,net228);
INTERCONNECT Split_269_n659_AND2T_62_n86(net229_c1,net229);
INTERCONNECT Split_277_n667_Split_278_n668(net230_c1,net230);
INTERCONNECT Split_285_n675_DFFT_128__FPB_n518(net231_c1,net231);
INTERCONNECT Split_293_n683_NOTT_18_n42(net232_c1,net232);
INTERCONNECT Split_301_n691_AND2T_93_n120(net233_c1,net233);
INTERCONNECT Split_278_n668_AND2T_22_n46(net234_c1,net234);
INTERCONNECT Split_286_n676_Split_287_n677(net235_c1,net235);
INTERCONNECT Split_294_n684_DFFT_136__FPB_n526(net236_c1,net236);
INTERCONNECT Split_302_n692_Split_303_n693(net237_c1,net237);
INTERCONNECT Split_279_n669_DFFT_131__FPB_n521(net238_c1,net238);
INTERCONNECT Split_287_n677_AND2T_31_n55(net239_c1,net239);
INTERCONNECT Split_295_n685_Split_296_n686(net240_c1,net240);
INTERCONNECT Split_303_n693_NOTT_10_n34(net241_c1,net241);
INTERCONNECT Split_288_n678_AND2T_58_n82(net242_c1,net242);
INTERCONNECT Split_296_n686_AND2T_70_n94(net243_c1,net243);
INTERCONNECT Split_304_n694_DFFT_135__FPB_n525(net244_c1,net244);
INTERCONNECT Split_289_n679_Split_290_n680(net245_c1,net245);
INTERCONNECT Split_297_n687_DFFT_185__FPB_n575(net246_c1,net246);
INTERCONNECT Split_305_n695_Split_306_n696(net247_c1,net247);
INTERCONNECT Split_298_n688_DFFT_119__FPB_n509(net248_c1,net248);
INTERCONNECT Split_306_n696_AND2T_14_n38(net249_c1,net249);
INTERCONNECT Split_299_n689_NOTT_8_n32(net250_c1,net250);
INTERCONNECT Split_307_n697_DFFT_117__FPB_n507(net251_c1,net251);
INTERCONNECT Split_308_n698_Split_309_n699(net252_c1,net252);
INTERCONNECT Split_309_n699_NOTT_12_n36(net253_c1,net253);
INTERCONNECT DFFT_100__PIPL_n136_DFFT_203__FPB_n593(net254_c1,net254);
INTERCONNECT DFFT_101__PIPL_n137_DFFT_210__FPB_n600(net255_c1,net255);
INTERCONNECT DFFT_102__PIPL_n138_DFFT_217__FPB_n607(net256_c1,net256);
INTERCONNECT DFFT_103__PIPL_n139_DFFT_224__FPB_n614(net257_c1,net257);
INTERCONNECT DFFT_110__FBL_n500_Split_305_n695(net258_c1,net258);
INTERCONNECT DFFT_111__FBL_n501_Split_308_n698(net259_c1,net259);
INTERCONNECT DFFT_104__FBL_n494_Split_298_n688(net260_c1,net260);
INTERCONNECT DFFT_105__FBL_n495_Split_300_n690(net261_c1,net261);
INTERCONNECT DFFT_106__FBL_n496_DFFT_202__FPB_n592(net262_c1,net262);
INTERCONNECT DFFT_107__FBL_n497_Split_301_n691(net263_c1,net263);
INTERCONNECT DFFT_108__FBL_n498_Split_302_n692(net264_c1,net264);
INTERCONNECT DFFT_109__FBL_n499_Split_HOLD_568(net265_c1,net265);
INTERCONNECT DFFT_98__FPB_n134_Split_292_n682(net266_c1,net266);
INTERCONNECT DFFT_99__FPB_n135_Split_295_n685(net267_c1,net267);
INTERCONNECT DFFT_112__FPB_n502_DFFT_106__FBL_n496(net268_c1,net268);
INTERCONNECT DFFT_120__FPB_n510_OR2T_27_n51(net269_c1,net269);
INTERCONNECT DFFT_113__FPB_n503_DFFT_107__FBL_n497(net270_c1,net270);
INTERCONNECT DFFT_121__FPB_n511_OR2T_28_n52(net271_c1,net271);
INTERCONNECT DFFT_210__FPB_n600_DFFT_211__FPB_n601(net272_c1,net272);
INTERCONNECT DFFT_122__FPB_n512_Split_HOLD_571(net273_c1,net273);
INTERCONNECT DFFT_114__FPB_n504_DFFT_109__FBL_n499(net274_c1,net274);
INTERCONNECT DFFT_130__FPB_n520_OR2T_34_n58(net275_c1,net275);
INTERCONNECT DFFT_211__FPB_n601_DFFT_212__FPB_n602(net276_c1,net276);
INTERCONNECT DFFT_123__FPB_n513_DFFT_124__FPB_n514(net277_c1,net277);
INTERCONNECT DFFT_115__FPB_n505_DFFT_110__FBL_n500(net278_c1,net278);
INTERCONNECT DFFT_131__FPB_n521_AND2T_36_n60(net279_c1,net279);
INTERCONNECT DFFT_220__FPB_n610_DFFT_221__FPB_n611(net280_c1,net280);
INTERCONNECT DFFT_212__FPB_n602_DFFT_213__FPB_n603(net281_c1,net281);
INTERCONNECT DFFT_132__FPB_n522_DFFT_133__FPB_n523(net282_c1,net282);
INTERCONNECT DFFT_124__FPB_n514_Split_HOLD_569(net283_c1,net283);
INTERCONNECT DFFT_116__FPB_n506_DFFT_111__FBL_n501(net284_c1,net284);
INTERCONNECT DFFT_140__FPB_n530_XOR2T_48_n72(net285_c1,net285);
INTERCONNECT DFFT_221__FPB_n611_DFFT_222__FPB_n612(net286_c1,net286);
INTERCONNECT DFFT_213__FPB_n603_Split_HOLD_567(net287_c1,net287);
INTERCONNECT DFFT_141__FPB_n531_OR2T_49_n73(net288_c1,net288);
INTERCONNECT DFFT_133__FPB_n523_OR2T_37_n61(net289_c1,net289);
INTERCONNECT DFFT_125__FPB_n515_AND2T_29_n53(net290_c1,net290);
INTERCONNECT DFFT_117__FPB_n507_AND2T_15_n39(net291_c1,net291);
INTERCONNECT DFFT_222__FPB_n612_DFFT_223_state_obs2(net292_c1,net292);
INTERCONNECT DFFT_214__FPB_n604_DFFT_215__FPB_n605(net293_c1,net293);
INTERCONNECT DFFT_150__FPB_n540_AND2T_53_n77(net294_c1,net294);
INTERCONNECT DFFT_142__FPB_n532_OR2T_50_n74(net295_c1,net295);
INTERCONNECT DFFT_134__FPB_n524_OR2T_38_n62(net296_c1,net296);
INTERCONNECT DFFT_126__FPB_n516_AND2T_30_n54(net297_c1,net297);
INTERCONNECT DFFT_118__FPB_n508_OR2T_16_n40(net298_c1,net298);
INTERCONNECT DFFT_215__FPB_n605_DFFT_216_state_obs1(net299_c1,net299);
INTERCONNECT DFFT_151__FPB_n541_OR2T_55_n79(net300_c1,net300);
INTERCONNECT DFFT_143__FPB_n533_OR2T_52_n76(net301_c1,net301);
INTERCONNECT DFFT_135__FPB_n525_AND2T_40_n64(net302_c1,net302);
INTERCONNECT DFFT_127__FPB_n517_AND2T_32_n56(net303_c1,net303);
INTERCONNECT DFFT_119__FPB_n509_AND2T_25_n49(net304_c1,net304);
INTERCONNECT DFFT_224__FPB_n614_DFFT_225__FPB_n615(net305_c1,net305);
INTERCONNECT DFFT_152__FPB_n542_DFFT_153__FPB_n543(net306_c1,net306);
INTERCONNECT DFFT_144__FPB_n534_DFFT_145__FPB_n535(net307_c1,net307);
INTERCONNECT DFFT_136__FPB_n526_Split_HOLD_566(net308_c1,net308);
INTERCONNECT DFFT_128__FPB_n518_DFFT_129__FPB_n519(net309_c1,net309);
INTERCONNECT DFFT_160__FPB_n550_AND2T_62_n86(net310_c1,net310);
INTERCONNECT DFFT_225__FPB_n615_DFFT_226__FPB_n616(net311_c1,net311);
INTERCONNECT DFFT_217__FPB_n607_DFFT_218__FPB_n608(net312_c1,net312);
INTERCONNECT DFFT_153__FPB_n543_DFFT_154__FPB_n544(net313_c1,net313);
INTERCONNECT DFFT_145__FPB_n535_DFFT_146__FPB_n536(net314_c1,net314);
INTERCONNECT DFFT_129__FPB_n519_DFFT_130__FPB_n520(net315_c1,net315);
INTERCONNECT DFFT_161__FPB_n551_AND2T_63_n87(net316_c1,net316);
INTERCONNECT DFFT_137__FPB_n527_AND2T_42_n66(net317_c1,net317);
INTERCONNECT DFFT_226__FPB_n616_DFFT_227__FPB_n617(net318_c1,net318);
INTERCONNECT DFFT_218__FPB_n608_DFFT_219__FPB_n609(net319_c1,net319);
INTERCONNECT DFFT_170__FPB_n560_DFFT_171__FPB_n561(net320_c1,net320);
INTERCONNECT DFFT_154__FPB_n544_DFFT_155__FPB_n545(net321_c1,net321);
INTERCONNECT DFFT_146__FPB_n536_DFFT_147__FPB_n537(net322_c1,net322);
INTERCONNECT DFFT_162__FPB_n552_OR2T_65_n89(net323_c1,net323);
INTERCONNECT DFFT_138__FPB_n528_AND2T_43_n67(net324_c1,net324);
INTERCONNECT DFFT_227__FPB_n617_DFFT_228__FPB_n618(net325_c1,net325);
INTERCONNECT DFFT_219__FPB_n609_DFFT_220__FPB_n610(net326_c1,net326);
INTERCONNECT DFFT_155__FPB_n545_DFFT_156__FPB_n546(net327_c1,net327);
INTERCONNECT DFFT_147__FPB_n537_DFFT_148__FPB_n538(net328_c1,net328);
INTERCONNECT DFFT_171__FPB_n561_AND2T_69_n93(net329_c1,net329);
INTERCONNECT DFFT_163__FPB_n553_OR2T_66_n90(net330_c1,net330);
INTERCONNECT DFFT_139__FPB_n529_AND2T_45_n69(net331_c1,net331);
INTERCONNECT DFFT_228__FPB_n618_DFFT_229_state_obs3(net332_c1,net332);
INTERCONNECT DFFT_180__FPB_n570_DFFT_181__FPB_n571(net333_c1,net333);
INTERCONNECT DFFT_148__FPB_n538_DFFT_149__FPB_n539(net334_c1,net334);
INTERCONNECT DFFT_172__FPB_n562_AND2T_70_n94(net335_c1,net335);
INTERCONNECT DFFT_164__FPB_n554_OR2T_67_n91(net336_c1,net336);
INTERCONNECT DFFT_156__FPB_n546_AND2T_56_n80(net337_c1,net337);
INTERCONNECT DFFT_181__FPB_n571_DFFT_182__FPB_n572(net338_c1,net338);
INTERCONNECT DFFT_165__FPB_n555_DFFT_166__FPB_n556(net339_c1,net339);
INTERCONNECT DFFT_157__FPB_n547_DFFT_158__FPB_n548(net340_c1,net340);
INTERCONNECT DFFT_149__FPB_n539_DFFT_150__FPB_n540(net341_c1,net341);
INTERCONNECT DFFT_173__FPB_n563_AND2T_74_n98(net342_c1,net342);
INTERCONNECT DFFT_190__FPB_n580_DFFT_191__FPB_n581(net343_c1,net343);
INTERCONNECT DFFT_182__FPB_n572_DFFT_183__FPB_n573(net344_c1,net344);
INTERCONNECT DFFT_174__FPB_n564_DFFT_175__FPB_n565(net345_c1,net345);
INTERCONNECT DFFT_166__FPB_n556_DFFT_167__FPB_n557(net346_c1,net346);
INTERCONNECT DFFT_158__FPB_n548_DFFT_159__FPB_n549(net347_c1,net347);
INTERCONNECT DFFT_183__FPB_n573_DFFT_184__FPB_n574(net348_c1,net348);
INTERCONNECT DFFT_167__FPB_n557_DFFT_168__FPB_n558(net349_c1,net349);
INTERCONNECT DFFT_191__FPB_n581_AND2T_85_n109(net350_c1,net350);
INTERCONNECT DFFT_175__FPB_n565_AND2T_76_n100(net351_c1,net351);
INTERCONNECT DFFT_159__FPB_n549_AND2T_60_n84(net352_c1,net352);
INTERCONNECT DFFT_168__FPB_n558_DFFT_169__FPB_n559(net353_c1,net353);
INTERCONNECT DFFT_200__FPB_n590_AND2T_92_n116(net354_c1,net354);
INTERCONNECT DFFT_192__FPB_n582_AND2T_86_n110(net355_c1,net355);
INTERCONNECT DFFT_184__FPB_n574_AND2T_82_n106(net356_c1,net356);
INTERCONNECT DFFT_176__FPB_n566_AND2T_77_n101(net357_c1,net357);
INTERCONNECT DFFT_185__FPB_n575_DFFT_186__FPB_n576(net358_c1,net358);
INTERCONNECT DFFT_169__FPB_n559_DFFT_170__FPB_n560(net359_c1,net359);
INTERCONNECT DFFT_201__FPB_n591_AND2T_94_n121(net360_c1,net360);
INTERCONNECT DFFT_193__FPB_n583_OR2T_90_n114(net361_c1,net361);
INTERCONNECT DFFT_177__FPB_n567_AND2T_78_n102(net362_c1,net362);
INTERCONNECT DFFT_186__FPB_n576_DFFT_187__FPB_n577(net363_c1,net363);
INTERCONNECT DFFT_202__FPB_n592_AND2T_96_n123(net364_c1,net364);
INTERCONNECT DFFT_194__FPB_n584_OR2T_91_n115(net365_c1,net365);
INTERCONNECT DFFT_178__FPB_n568_OR2T_81_n105(net366_c1,net366);
INTERCONNECT DFFT_203__FPB_n593_Split_HOLD_570(net367_c1,net367);
INTERCONNECT DFFT_195__FPB_n585_DFFT_196__FPB_n586(net368_c1,net368);
INTERCONNECT DFFT_179__FPB_n569_DFFT_180__FPB_n570(net369_c1,net369);
INTERCONNECT DFFT_187__FPB_n577_AND2T_83_n107(net370_c1,net370);
INTERCONNECT DFFT_204__FPB_n594_DFFT_205__FPB_n595(net371_c1,net371);
INTERCONNECT DFFT_196__FPB_n586_DFFT_197__FPB_n587(net372_c1,net372);
INTERCONNECT DFFT_188__FPB_n578_DFFT_189__FPB_n579(net373_c1,net373);
INTERCONNECT DFFT_205__FPB_n595_DFFT_206__FPB_n596(net374_c1,net374);
INTERCONNECT DFFT_197__FPB_n587_DFFT_198__FPB_n588(net375_c1,net375);
INTERCONNECT DFFT_189__FPB_n579_AND2T_84_n108(net376_c1,net376);
INTERCONNECT DFFT_206__FPB_n596_DFFT_207__FPB_n597(net377_c1,net377);
INTERCONNECT DFFT_198__FPB_n588_DFFT_199__FPB_n589(net378_c1,net378);
INTERCONNECT DFFT_207__FPB_n597_DFFT_208__FPB_n598(net379_c1,net379);
INTERCONNECT DFFT_199__FPB_n589_DFFT_200__FPB_n590(net380_c1,net380);
INTERCONNECT DFFT_208__FPB_n598_DFFT_209_state_obs0(net381_c1,net381);
INTERCONNECT DFFT_209_state_obs0_state_obs0_Pad(net382_c1,state_obs0_Pad);
INTERCONNECT DFFT_216_state_obs1_state_obs1_Pad(net383_c1,state_obs1_Pad);
INTERCONNECT DFFT_223_state_obs2_state_obs2_Pad(net384_c1,state_obs2_Pad);
INTERCONNECT DFFT_229_state_obs3_state_obs3_Pad(net385_c1,state_obs3_Pad);
INTERCONNECT SplitCLK_0_477_SplitCLK_0_332(net386_c1,net386);
INTERCONNECT SplitCLK_0_477_SplitCLK_2_442(net387_c1,net387);
INTERCONNECT SplitCLK_2_476_DFFT_98__FPB_n134(net388_c1,net388);
INTERCONNECT SplitCLK_2_475_DFFT_197__FPB_n587(net389_c1,net389);
INTERCONNECT SplitCLK_2_474_DFFT_185__FPB_n575(net390_c1,net390);
INTERCONNECT SplitCLK_2_473_DFFT_168__FPB_n558(net391_c1,net391);
INTERCONNECT SplitCLK_2_472_DFFT_159__FPB_n549(net392_c1,net392);
INTERCONNECT SplitCLK_2_471_DFFT_183__FPB_n573(net393_c1,net393);
INTERCONNECT SplitCLK_2_470_DFFT_174__FPB_n564(net394_c1,net394);
INTERCONNECT SplitCLK_2_469_DFFT_148__FPB_n538(net395_c1,net395);
INTERCONNECT SplitCLK_2_468_DFFT_146__FPB_n536(net396_c1,net396);
INTERCONNECT SplitCLK_2_467_DFFT_217__FPB_n607(net397_c1,net397);
INTERCONNECT SplitCLK_2_466_DFFT_128__FPB_n518(net398_c1,net398);
INTERCONNECT SplitCLK_2_465_DFFT_136__FPB_n526(net399_c1,net399);
INTERCONNECT SplitCLK_2_464_DFFT_143__FPB_n533(net400_c1,net400);
INTERCONNECT SplitCLK_2_463_DFFT_141__FPB_n531(net401_c1,net401);
INTERCONNECT SplitCLK_2_462_DFFT_116__FPB_n506(net402_c1,net402);
INTERCONNECT SplitCLK_2_461_DFFT_124__FPB_n514(net403_c1,net403);
INTERCONNECT SplitCLK_2_460_DFFT_107__FBL_n497(net404_c1,net404);
INTERCONNECT SplitCLK_4_459_DFFT_104__FBL_n494(net405_c1,net405);
INTERCONNECT SplitCLK_4_458_AND2T_96_n123(net406_c1,net406);
INTERCONNECT SplitCLK_2_457_AND2T_78_n102(net407_c1,net407);
INTERCONNECT SplitCLK_2_456_AND2T_85_n109(net408_c1,net408);
INTERCONNECT SplitCLK_2_455_NOTT_23_n47(net409_c1,net409);
INTERCONNECT SplitCLK_2_454_NOTT_13_n37(net410_c1,net410);
INTERCONNECT SplitCLK_2_453_NOTT_11_n35(net411_c1,net411);
INTERCONNECT SplitCLK_2_452_OR2T_75_n99(net412_c1,net412);
INTERCONNECT SplitCLK_2_451_OR2T_66_n90(net413_c1,net413);
INTERCONNECT SplitCLK_2_450_OR2T_46_n70(net414_c1,net414);
INTERCONNECT SplitCLK_2_449_AND2T_57_n81(net415_c1,net415);
INTERCONNECT SplitCLK_2_448_AND2T_56_n80(net416_c1,net416);
INTERCONNECT SplitCLK_2_447_AND2T_53_n77(net417_c1,net417);
INTERCONNECT SplitCLK_4_446_AND2T_43_n67(net418_c1,net418);
INTERCONNECT SplitCLK_2_445_AND2T_25_n49(net419_c1,net419);
INTERCONNECT SplitCLK_2_444_AND2T_31_n55(net420_c1,net420);
INTERCONNECT SplitCLK_2_443_NOTT_9_n33(net421_c1,net421);
INTERCONNECT SplitCLK_2_442_SplitCLK_6_387(net422_c1,net422);
INTERCONNECT SplitCLK_2_442_SplitCLK_4_441(net423_c1,net423);
INTERCONNECT SplitCLK_4_441_SplitCLK_0_414(net424_c1,net424);
INTERCONNECT SplitCLK_4_441_SplitCLK_2_440(net425_c1,net425);
INTERCONNECT SplitCLK_2_440_SplitCLK_6_427(net426_c1,net426);
INTERCONNECT SplitCLK_2_440_SplitCLK_4_439(net427_c1,net427);
INTERCONNECT SplitCLK_4_439_SplitCLK_0_433(net428_c1,net428);
INTERCONNECT SplitCLK_4_439_SplitCLK_2_438(net429_c1,net429);
INTERCONNECT SplitCLK_2_438_SplitCLK_2_435(net430_c1,net430);
INTERCONNECT SplitCLK_2_438_SplitCLK_2_437(net431_c1,net431);
INTERCONNECT SplitCLK_2_437_SplitCLK_2_469(net432_c1,net432);
INTERCONNECT SplitCLK_2_437_SplitCLK_4_436(net433_c1,net433);
INTERCONNECT SplitCLK_4_436_DFFT_147__FPB_n537(net434_c1,net434);
INTERCONNECT SplitCLK_4_436_DFFT_149__FPB_n539(net435_c1,net435);
INTERCONNECT SplitCLK_2_435_SplitCLK_2_461(net436_c1,net436);
INTERCONNECT SplitCLK_2_435_SplitCLK_4_434(net437_c1,net437);
INTERCONNECT SplitCLK_4_434_DFFT_150__FPB_n540(net438_c1,net438);
INTERCONNECT SplitCLK_4_434_DFFT_152__FPB_n542(net439_c1,net439);
INTERCONNECT SplitCLK_0_433_SplitCLK_0_430(net440_c1,net440);
INTERCONNECT SplitCLK_0_433_SplitCLK_4_432(net441_c1,net441);
INTERCONNECT SplitCLK_4_432_SplitCLK_2_468(net442_c1,net442);
INTERCONNECT SplitCLK_4_432_SplitCLK_4_431(net443_c1,net443);
INTERCONNECT SplitCLK_4_431_DFFT_144__FPB_n534(net444_c1,net444);
INTERCONNECT SplitCLK_4_431_DFFT_145__FPB_n535(net445_c1,net445);
INTERCONNECT SplitCLK_0_430_SplitCLK_4_428(net446_c1,net446);
INTERCONNECT SplitCLK_0_430_SplitCLK_4_429(net447_c1,net447);
INTERCONNECT SplitCLK_4_429_DFFT_153__FPB_n543(net448_c1,net448);
INTERCONNECT SplitCLK_4_429_NOTT_95_n122(net449_c1,net449);
INTERCONNECT SplitCLK_4_428_DFFT_122__FPB_n512(net450_c1,net450);
INTERCONNECT SplitCLK_4_428_DFFT_154__FPB_n544(net451_c1,net451);
INTERCONNECT SplitCLK_6_427_SplitCLK_0_420(net452_c1,net452);
INTERCONNECT SplitCLK_6_427_SplitCLK_2_426(net453_c1,net453);
INTERCONNECT SplitCLK_2_426_SplitCLK_2_423(net454_c1,net454);
INTERCONNECT SplitCLK_2_426_SplitCLK_4_425(net455_c1,net455);
INTERCONNECT SplitCLK_4_425_SplitCLK_2_447(net456_c1,net456);
INTERCONNECT SplitCLK_4_425_SplitCLK_4_424(net457_c1,net457);
INTERCONNECT SplitCLK_4_424_DFFT_123__FPB_n513(net458_c1,net458);
INTERCONNECT SplitCLK_4_424_DFFT_125__FPB_n515(net459_c1,net459);
INTERCONNECT SplitCLK_2_423_SplitCLK_4_421(net460_c1,net460);
INTERCONNECT SplitCLK_2_423_SplitCLK_4_422(net461_c1,net461);
INTERCONNECT SplitCLK_4_422_OR2T_51_n75(net462_c1,net462);
INTERCONNECT SplitCLK_4_422_DFFT_138__FPB_n528(net463_c1,net463);
INTERCONNECT SplitCLK_4_421_OR2T_50_n74(net464_c1,net464);
INTERCONNECT SplitCLK_4_421_OR2T_52_n76(net465_c1,net465);
INTERCONNECT SplitCLK_0_420_SplitCLK_4_417(net466_c1,net466);
INTERCONNECT SplitCLK_0_420_SplitCLK_4_419(net467_c1,net467);
INTERCONNECT SplitCLK_4_419_SplitCLK_2_464(net468_c1,net468);
INTERCONNECT SplitCLK_4_419_SplitCLK_4_418(net469_c1,net469);
INTERCONNECT SplitCLK_4_418_AND2T_29_n53(net470_c1,net470);
INTERCONNECT SplitCLK_4_418_DFFT_137__FPB_n527(net471_c1,net471);
INTERCONNECT SplitCLK_4_417_SplitCLK_4_415(net472_c1,net472);
INTERCONNECT SplitCLK_4_417_SplitCLK_4_416(net473_c1,net473);
INTERCONNECT SplitCLK_4_416_AND2T_42_n66(net474_c1,net474);
INTERCONNECT SplitCLK_4_416_DFFT_142__FPB_n532(net475_c1,net475);
INTERCONNECT SplitCLK_4_415_AND2T_39_n63(net476_c1,net476);
INTERCONNECT SplitCLK_4_415_OR2T_37_n61(net477_c1,net477);
INTERCONNECT SplitCLK_0_414_SplitCLK_6_400(net478_c1,net478);
INTERCONNECT SplitCLK_0_414_SplitCLK_4_413(net479_c1,net479);
INTERCONNECT SplitCLK_4_413_SplitCLK_4_406(net480_c1,net480);
INTERCONNECT SplitCLK_4_413_SplitCLK_6_412(net481_c1,net481);
INTERCONNECT SplitCLK_6_412_SplitCLK_4_409(net482_c1,net482);
INTERCONNECT SplitCLK_6_412_SplitCLK_2_411(net483_c1,net483);
INTERCONNECT SplitCLK_2_411_SplitCLK_2_476(net484_c1,net484);
INTERCONNECT SplitCLK_2_411_SplitCLK_4_410(net485_c1,net485);
INTERCONNECT SplitCLK_4_410_DFFT_165__FPB_n555(net486_c1,net486);
INTERCONNECT SplitCLK_4_410_DFFT_166__FPB_n556(net487_c1,net487);
INTERCONNECT SplitCLK_4_409_SplitCLK_0_407(net488_c1,net488);
INTERCONNECT SplitCLK_4_409_SplitCLK_4_408(net489_c1,net489);
INTERCONNECT SplitCLK_4_408_DFFT_170__FPB_n560(net490_c1,net490);
INTERCONNECT SplitCLK_4_408_DFFT_156__FPB_n546(net491_c1,net491);
INTERCONNECT SplitCLK_0_407_AND2T_69_n93(net492_c1,net492);
INTERCONNECT SplitCLK_0_407_DFFT_169__FPB_n559(net493_c1,net493);
INTERCONNECT SplitCLK_4_406_SplitCLK_6_403(net494_c1,net494);
INTERCONNECT SplitCLK_4_406_SplitCLK_4_405(net495_c1,net495);
INTERCONNECT SplitCLK_4_405_SplitCLK_2_473(net496_c1,net496);
INTERCONNECT SplitCLK_4_405_SplitCLK_4_404(net497_c1,net497);
INTERCONNECT SplitCLK_4_404_DFFT_181__FPB_n571(net498_c1,net498);
INTERCONNECT SplitCLK_4_404_DFFT_167__FPB_n557(net499_c1,net499);
INTERCONNECT SplitCLK_6_403_SplitCLK_4_401(net500_c1,net500);
INTERCONNECT SplitCLK_6_403_SplitCLK_4_402(net501_c1,net501);
INTERCONNECT SplitCLK_4_402_OR2T_68_n92(net502_c1,net502);
INTERCONNECT SplitCLK_4_402_DFFT_171__FPB_n561(net503_c1,net503);
INTERCONNECT SplitCLK_4_401_DFFT_157__FPB_n547(net504_c1,net504);
INTERCONNECT SplitCLK_4_401_DFFT_158__FPB_n548(net505_c1,net505);
INTERCONNECT SplitCLK_6_400_SplitCLK_0_393(net506_c1,net506);
INTERCONNECT SplitCLK_6_400_SplitCLK_2_399(net507_c1,net507);
INTERCONNECT SplitCLK_2_399_SplitCLK_2_396(net508_c1,net508);
INTERCONNECT SplitCLK_2_399_SplitCLK_2_398(net509_c1,net509);
INTERCONNECT SplitCLK_2_398_SplitCLK_2_465(net510_c1,net510);
INTERCONNECT SplitCLK_2_398_SplitCLK_4_397(net511_c1,net511);
INTERCONNECT SplitCLK_4_397_DFFT_108__FBL_n498(net512_c1,net512);
INTERCONNECT SplitCLK_4_397_DFFT_155__FPB_n545(net513_c1,net513);
INTERCONNECT SplitCLK_2_396_SplitCLK_4_394(net514_c1,net514);
INTERCONNECT SplitCLK_2_396_SplitCLK_4_395(net515_c1,net515);
INTERCONNECT SplitCLK_4_395_DFFT_132__FPB_n522(net516_c1,net516);
INTERCONNECT SplitCLK_4_395_DFFT_133__FPB_n523(net517_c1,net517);
INTERCONNECT SplitCLK_4_394_OR2T_54_n78(net518_c1,net518);
INTERCONNECT SplitCLK_4_394_DFFT_151__FPB_n541(net519_c1,net519);
INTERCONNECT SplitCLK_0_393_SplitCLK_6_390(net520_c1,net520);
INTERCONNECT SplitCLK_0_393_SplitCLK_4_392(net521_c1,net521);
INTERCONNECT SplitCLK_4_392_SplitCLK_2_448(net522_c1,net522);
INTERCONNECT SplitCLK_4_392_SplitCLK_4_391(net523_c1,net523);
INTERCONNECT SplitCLK_4_391_DFFT_130__FPB_n520(net524_c1,net524);
INTERCONNECT SplitCLK_4_391_DFFT_129__FPB_n519(net525_c1,net525);
INTERCONNECT SplitCLK_6_390_SplitCLK_4_388(net526_c1,net526);
INTERCONNECT SplitCLK_6_390_SplitCLK_4_389(net527_c1,net527);
INTERCONNECT SplitCLK_4_389_OR2T_34_n58(net528_c1,net528);
INTERCONNECT SplitCLK_4_389_OR2T_55_n79(net529_c1,net529);
INTERCONNECT SplitCLK_4_388_OR2T_64_n88(net530_c1,net530);
INTERCONNECT SplitCLK_4_388_NOTT_18_n42(net531_c1,net531);
INTERCONNECT SplitCLK_6_387_SplitCLK_6_359(net532_c1,net532);
INTERCONNECT SplitCLK_6_387_SplitCLK_2_386(net533_c1,net533);
INTERCONNECT SplitCLK_2_386_SplitCLK_6_372(net534_c1,net534);
INTERCONNECT SplitCLK_2_386_SplitCLK_4_385(net535_c1,net535);
INTERCONNECT SplitCLK_4_385_SplitCLK_4_378(net536_c1,net536);
INTERCONNECT SplitCLK_4_385_SplitCLK_2_384(net537_c1,net537);
INTERCONNECT SplitCLK_2_384_SplitCLK_6_381(net538_c1,net538);
INTERCONNECT SplitCLK_2_384_SplitCLK_4_383(net539_c1,net539);
INTERCONNECT SplitCLK_4_383_SplitCLK_4_459(net540_c1,net540);
INTERCONNECT SplitCLK_4_383_SplitCLK_4_382(net541_c1,net541);
INTERCONNECT SplitCLK_4_382_AND2T_40_n64(net542_c1,net542);
INTERCONNECT SplitCLK_4_382_DFFT_135__FPB_n525(net543_c1,net543);
INTERCONNECT SplitCLK_6_381_SplitCLK_4_379(net544_c1,net544);
INTERCONNECT SplitCLK_6_381_SplitCLK_4_380(net545_c1,net545);
INTERCONNECT SplitCLK_4_380_NOTT_8_n32(net546_c1,net546);
INTERCONNECT SplitCLK_4_380_NOTT_12_n36(net547_c1,net547);
INTERCONNECT SplitCLK_4_379_AND2T_94_n121(net548_c1,net548);
INTERCONNECT SplitCLK_4_379_DFFT_119__FPB_n509(net549_c1,net549);
INTERCONNECT SplitCLK_4_378_SplitCLK_0_375(net550_c1,net550);
INTERCONNECT SplitCLK_4_378_SplitCLK_4_377(net551_c1,net551);
INTERCONNECT SplitCLK_4_377_SplitCLK_4_446(net552_c1,net552);
INTERCONNECT SplitCLK_4_377_SplitCLK_4_376(net553_c1,net553);
INTERCONNECT SplitCLK_4_376_OR2T_38_n62(net554_c1,net554);
INTERCONNECT SplitCLK_4_376_DFFT_134__FPB_n524(net555_c1,net555);
INTERCONNECT SplitCLK_0_375_SplitCLK_4_373(net556_c1,net556);
INTERCONNECT SplitCLK_0_375_SplitCLK_0_374(net557_c1,net557);
INTERCONNECT SplitCLK_0_374_AND2T_21_n45(net558_c1,net558);
INTERCONNECT SplitCLK_0_374_DFFT_201__FPB_n591(net559_c1,net559);
INTERCONNECT SplitCLK_4_373_AND2T_35_n59(net560_c1,net560);
INTERCONNECT SplitCLK_4_373_NOTT_10_n34(net561_c1,net561);
INTERCONNECT SplitCLK_6_372_SplitCLK_4_365(net562_c1,net562);
INTERCONNECT SplitCLK_6_372_SplitCLK_2_371(net563_c1,net563);
INTERCONNECT SplitCLK_2_371_SplitCLK_4_368(net564_c1,net564);
INTERCONNECT SplitCLK_2_371_SplitCLK_2_370(net565_c1,net565);
INTERCONNECT SplitCLK_2_370_SplitCLK_2_462(net566_c1,net566);
INTERCONNECT SplitCLK_2_370_SplitCLK_4_369(net567_c1,net567);
INTERCONNECT SplitCLK_4_369_DFFT_111__FBL_n501(net568_c1,net568);
INTERCONNECT SplitCLK_4_369_DFFT_204__FPB_n594(net569_c1,net569);
INTERCONNECT SplitCLK_4_368_SplitCLK_4_366(net570_c1,net570);
INTERCONNECT SplitCLK_4_368_SplitCLK_4_367(net571_c1,net571);
INTERCONNECT SplitCLK_4_367_DFFT_209_state_obs0(net572_c1,net572);
INTERCONNECT SplitCLK_4_367_DFFT_203__FPB_n593(net573_c1,net573);
INTERCONNECT SplitCLK_4_366_DFFT_100__PIPL_n136(net574_c1,net574);
INTERCONNECT SplitCLK_4_366_DFFT_208__FPB_n598(net575_c1,net575);
INTERCONNECT SplitCLK_4_365_SplitCLK_0_362(net576_c1,net576);
INTERCONNECT SplitCLK_4_365_SplitCLK_0_364(net577_c1,net577);
INTERCONNECT SplitCLK_0_364_SplitCLK_2_443(net578_c1,net578);
INTERCONNECT SplitCLK_0_364_SplitCLK_4_363(net579_c1,net579);
INTERCONNECT SplitCLK_4_363_DFFT_106__FBL_n496(net580_c1,net580);
INTERCONNECT SplitCLK_4_363_DFFT_202__FPB_n592(net581_c1,net581);
INTERCONNECT SplitCLK_0_362_SplitCLK_4_360(net582_c1,net582);
INTERCONNECT SplitCLK_0_362_SplitCLK_0_361(net583_c1,net583);
INTERCONNECT SplitCLK_0_361_DFFT_206__FPB_n596(net584_c1,net584);
INTERCONNECT SplitCLK_0_361_DFFT_207__FPB_n597(net585_c1,net585);
INTERCONNECT SplitCLK_4_360_DFFT_101__PIPL_n137(net586_c1,net586);
INTERCONNECT SplitCLK_4_360_DFFT_205__FPB_n595(net587_c1,net587);
INTERCONNECT SplitCLK_6_359_SplitCLK_6_345(net588_c1,net588);
INTERCONNECT SplitCLK_6_359_SplitCLK_4_358(net589_c1,net589);
INTERCONNECT SplitCLK_4_358_SplitCLK_4_351(net590_c1,net590);
INTERCONNECT SplitCLK_4_358_SplitCLK_2_357(net591_c1,net591);
INTERCONNECT SplitCLK_2_357_SplitCLK_6_354(net592_c1,net592);
INTERCONNECT SplitCLK_2_357_SplitCLK_4_356(net593_c1,net593);
INTERCONNECT SplitCLK_4_356_SplitCLK_2_445(net594_c1,net594);
INTERCONNECT SplitCLK_4_356_SplitCLK_4_355(net595_c1,net595);
INTERCONNECT SplitCLK_4_355_AND2T_45_n69(net596_c1,net596);
INTERCONNECT SplitCLK_4_355_OR2T_87_n111(net597_c1,net597);
INTERCONNECT SplitCLK_6_354_SplitCLK_4_352(net598_c1,net598);
INTERCONNECT SplitCLK_6_354_SplitCLK_0_353(net599_c1,net599);
INTERCONNECT SplitCLK_0_353_AND2T_19_n43(net600_c1,net600);
INTERCONNECT SplitCLK_0_353_AND2T_93_n120(net601_c1,net601);
INTERCONNECT SplitCLK_4_352_DFFT_118__FPB_n508(net602_c1,net602);
INTERCONNECT SplitCLK_4_352_DFFT_139__FPB_n529(net603_c1,net603);
INTERCONNECT SplitCLK_4_351_SplitCLK_0_348(net604_c1,net604);
INTERCONNECT SplitCLK_4_351_SplitCLK_2_350(net605_c1,net605);
INTERCONNECT SplitCLK_2_350_SplitCLK_2_463(net606_c1,net606);
INTERCONNECT SplitCLK_2_350_SplitCLK_4_349(net607_c1,net607);
INTERCONNECT SplitCLK_4_349_AND2T_47_n71(net608_c1,net608);
INTERCONNECT SplitCLK_4_349_OR2T_49_n73(net609_c1,net609);
INTERCONNECT SplitCLK_0_348_SplitCLK_4_346(net610_c1,net610);
INTERCONNECT SplitCLK_0_348_SplitCLK_0_347(net611_c1,net611);
INTERCONNECT SplitCLK_0_347_OR2T_28_n52(net612_c1,net612);
INTERCONNECT SplitCLK_0_347_DFFT_131__FPB_n521(net613_c1,net613);
INTERCONNECT SplitCLK_4_346_AND2T_36_n60(net614_c1,net614);
INTERCONNECT SplitCLK_4_346_DFFT_121__FPB_n511(net615_c1,net615);
INTERCONNECT SplitCLK_6_345_SplitCLK_4_338(net616_c1,net616);
INTERCONNECT SplitCLK_6_345_SplitCLK_2_344(net617_c1,net617);
INTERCONNECT SplitCLK_2_344_SplitCLK_0_341(net618_c1,net618);
INTERCONNECT SplitCLK_2_344_SplitCLK_2_343(net619_c1,net619);
INTERCONNECT SplitCLK_2_343_SplitCLK_2_453(net620_c1,net620);
INTERCONNECT SplitCLK_2_343_SplitCLK_4_342(net621_c1,net621);
INTERCONNECT SplitCLK_4_342_DFFT_112__FPB_n502(net622_c1,net622);
INTERCONNECT SplitCLK_4_342_DFFT_210__FPB_n600(net623_c1,net623);
INTERCONNECT SplitCLK_0_341_SplitCLK_4_339(net624_c1,net624);
INTERCONNECT SplitCLK_0_341_SplitCLK_0_340(net625_c1,net625);
INTERCONNECT SplitCLK_0_340_DFFT_212__FPB_n602(net626_c1,net626);
INTERCONNECT SplitCLK_0_340_DFFT_216_state_obs1(net627_c1,net627);
INTERCONNECT SplitCLK_4_339_DFFT_211__FPB_n601(net628_c1,net628);
INTERCONNECT SplitCLK_4_339_DFFT_213__FPB_n603(net629_c1,net629);
INTERCONNECT SplitCLK_4_338_SplitCLK_0_335(net630_c1,net630);
INTERCONNECT SplitCLK_4_338_SplitCLK_6_337(net631_c1,net631);
INTERCONNECT SplitCLK_6_337_SplitCLK_4_458(net632_c1,net632);
INTERCONNECT SplitCLK_6_337_SplitCLK_4_336(net633_c1,net633);
INTERCONNECT SplitCLK_4_336_XOR2T_48_n72(net634_c1,net634);
INTERCONNECT SplitCLK_4_336_DFFT_114__FPB_n504(net635_c1,net635);
INTERCONNECT SplitCLK_0_335_SplitCLK_4_333(net636_c1,net636);
INTERCONNECT SplitCLK_0_335_SplitCLK_0_334(net637_c1,net637);
INTERCONNECT SplitCLK_0_334_DFFT_214__FPB_n604(net638_c1,net638);
INTERCONNECT SplitCLK_0_334_DFFT_215__FPB_n605(net639_c1,net639);
INTERCONNECT SplitCLK_4_333_DFFT_109__FBL_n499(net640_c1,net640);
INTERCONNECT SplitCLK_4_333_DFFT_223_state_obs2(net641_c1,net641);
INTERCONNECT SplitCLK_0_332_SplitCLK_6_277(net642_c1,net642);
INTERCONNECT SplitCLK_0_332_SplitCLK_4_331(net643_c1,net643);
INTERCONNECT SplitCLK_4_331_SplitCLK_0_304(net644_c1,net644);
INTERCONNECT SplitCLK_4_331_SplitCLK_2_330(net645_c1,net645);
INTERCONNECT SplitCLK_2_330_SplitCLK_6_317(net646_c1,net646);
INTERCONNECT SplitCLK_2_330_SplitCLK_4_329(net647_c1,net647);
INTERCONNECT SplitCLK_4_329_SplitCLK_0_323(net648_c1,net648);
INTERCONNECT SplitCLK_4_329_SplitCLK_6_328(net649_c1,net649);
INTERCONNECT SplitCLK_6_328_SplitCLK_2_325(net650_c1,net650);
INTERCONNECT SplitCLK_6_328_SplitCLK_4_327(net651_c1,net651);
INTERCONNECT SplitCLK_4_327_SplitCLK_2_472(net652_c1,net652);
INTERCONNECT SplitCLK_4_327_SplitCLK_4_326(net653_c1,net653);
INTERCONNECT SplitCLK_4_326_DFFT_180__FPB_n570(net654_c1,net654);
INTERCONNECT SplitCLK_4_326_DFFT_182__FPB_n572(net655_c1,net655);
INTERCONNECT SplitCLK_2_325_SplitCLK_2_466(net656_c1,net656);
INTERCONNECT SplitCLK_2_325_SplitCLK_4_324(net657_c1,net657);
INTERCONNECT SplitCLK_4_324_DFFT_99__FPB_n135(net658_c1,net658);
INTERCONNECT SplitCLK_4_324_OR2T_67_n91(net659_c1,net659);
INTERCONNECT SplitCLK_0_323_SplitCLK_6_320(net660_c1,net660);
INTERCONNECT SplitCLK_0_323_SplitCLK_4_322(net661_c1,net661);
INTERCONNECT SplitCLK_4_322_SplitCLK_2_471(net662_c1,net662);
INTERCONNECT SplitCLK_4_322_SplitCLK_4_321(net663_c1,net663);
INTERCONNECT SplitCLK_4_321_NOTT_17_n41(net664_c1,net664);
INTERCONNECT SplitCLK_4_321_DFFT_179__FPB_n569(net665_c1,net665);
INTERCONNECT SplitCLK_6_320_SplitCLK_4_318(net666_c1,net666);
INTERCONNECT SplitCLK_6_320_SplitCLK_4_319(net667_c1,net667);
INTERCONNECT SplitCLK_4_319_AND2T_60_n84(net668_c1,net668);
INTERCONNECT SplitCLK_4_319_DFFT_164__FPB_n554(net669_c1,net669);
INTERCONNECT SplitCLK_4_318_DFFT_184__FPB_n574(net670_c1,net670);
INTERCONNECT SplitCLK_4_318_DFFT_188__FPB_n578(net671_c1,net671);
INTERCONNECT SplitCLK_6_317_SplitCLK_4_310(net672_c1,net672);
INTERCONNECT SplitCLK_6_317_SplitCLK_2_316(net673_c1,net673);
INTERCONNECT SplitCLK_2_316_SplitCLK_6_313(net674_c1,net674);
INTERCONNECT SplitCLK_2_316_SplitCLK_4_315(net675_c1,net675);
INTERCONNECT SplitCLK_4_315_SplitCLK_2_451(net676_c1,net676);
INTERCONNECT SplitCLK_4_315_SplitCLK_4_314(net677_c1,net677);
INTERCONNECT SplitCLK_4_314_DFFT_105__FBL_n495(net678_c1,net678);
INTERCONNECT SplitCLK_4_314_DFFT_172__FPB_n562(net679_c1,net679);
INTERCONNECT SplitCLK_6_313_SplitCLK_4_311(net680_c1,net680);
INTERCONNECT SplitCLK_6_313_SplitCLK_0_312(net681_c1,net681);
INTERCONNECT SplitCLK_0_312_OR2T_65_n89(net682_c1,net682);
INTERCONNECT SplitCLK_0_312_DFFT_163__FPB_n553(net683_c1,net683);
INTERCONNECT SplitCLK_4_311_DFFT_162__FPB_n552(net684_c1,net684);
INTERCONNECT SplitCLK_4_311_DFFT_177__FPB_n567(net685_c1,net685);
INTERCONNECT SplitCLK_4_310_SplitCLK_0_307(net686_c1,net686);
INTERCONNECT SplitCLK_4_310_SplitCLK_2_309(net687_c1,net687);
INTERCONNECT SplitCLK_2_309_SplitCLK_2_457(net688_c1,net688);
INTERCONNECT SplitCLK_2_309_SplitCLK_4_308(net689_c1,net689);
INTERCONNECT SplitCLK_4_308_AND2T_70_n94(net690_c1,net690);
INTERCONNECT SplitCLK_4_308_DFFT_190__FPB_n580(net691_c1,net691);
INTERCONNECT SplitCLK_0_307_SplitCLK_4_305(net692_c1,net692);
INTERCONNECT SplitCLK_0_307_SplitCLK_0_306(net693_c1,net693);
INTERCONNECT SplitCLK_0_306_AND2T_82_n106(net694_c1,net694);
INTERCONNECT SplitCLK_0_306_OR2T_81_n105(net695_c1,net695);
INTERCONNECT SplitCLK_4_305_AND2T_71_n95(net696_c1,net696);
INTERCONNECT SplitCLK_4_305_OR2T_80_n104(net697_c1,net697);
INTERCONNECT SplitCLK_0_304_SplitCLK_6_290(net698_c1,net698);
INTERCONNECT SplitCLK_0_304_SplitCLK_4_303(net699_c1,net699);
INTERCONNECT SplitCLK_4_303_SplitCLK_0_296(net700_c1,net700);
INTERCONNECT SplitCLK_4_303_SplitCLK_2_302(net701_c1,net701);
INTERCONNECT SplitCLK_2_302_SplitCLK_4_299(net702_c1,net702);
INTERCONNECT SplitCLK_2_302_SplitCLK_4_301(net703_c1,net703);
INTERCONNECT SplitCLK_4_301_SplitCLK_2_474(net704_c1,net704);
INTERCONNECT SplitCLK_4_301_SplitCLK_4_300(net705_c1,net705);
INTERCONNECT SplitCLK_4_300_DFFT_195__FPB_n585(net706_c1,net706);
INTERCONNECT SplitCLK_4_300_DFFT_196__FPB_n586(net707_c1,net707);
INTERCONNECT SplitCLK_4_299_SplitCLK_4_297(net708_c1,net708);
INTERCONNECT SplitCLK_4_299_SplitCLK_4_298(net709_c1,net709);
INTERCONNECT SplitCLK_4_298_DFFT_186__FPB_n576(net710_c1,net710);
INTERCONNECT SplitCLK_4_298_DFFT_189__FPB_n579(net711_c1,net711);
INTERCONNECT SplitCLK_4_297_AND2T_83_n107(net712_c1,net712);
INTERCONNECT SplitCLK_4_297_DFFT_187__FPB_n577(net713_c1,net713);
INTERCONNECT SplitCLK_0_296_SplitCLK_4_293(net714_c1,net714);
INTERCONNECT SplitCLK_0_296_SplitCLK_4_295(net715_c1,net715);
INTERCONNECT SplitCLK_4_295_SplitCLK_2_475(net716_c1,net716);
INTERCONNECT SplitCLK_4_295_SplitCLK_4_294(net717_c1,net717);
INTERCONNECT SplitCLK_4_294_DFFT_200__FPB_n590(net718_c1,net718);
INTERCONNECT SplitCLK_4_294_DFFT_198__FPB_n588(net719_c1,net719);
INTERCONNECT SplitCLK_4_293_SplitCLK_4_291(net720_c1,net720);
INTERCONNECT SplitCLK_4_293_SplitCLK_4_292(net721_c1,net721);
INTERCONNECT SplitCLK_4_292_OR2T_91_n115(net722_c1,net722);
INTERCONNECT SplitCLK_4_292_DFFT_194__FPB_n584(net723_c1,net723);
INTERCONNECT SplitCLK_4_291_DFFT_199__FPB_n589(net724_c1,net724);
INTERCONNECT SplitCLK_4_291_AND2T_92_n116(net725_c1,net725);
INTERCONNECT SplitCLK_6_290_SplitCLK_4_283(net726_c1,net726);
INTERCONNECT SplitCLK_6_290_SplitCLK_2_289(net727_c1,net727);
INTERCONNECT SplitCLK_2_289_SplitCLK_6_286(net728_c1,net728);
INTERCONNECT SplitCLK_2_289_SplitCLK_4_288(net729_c1,net729);
INTERCONNECT SplitCLK_4_288_SplitCLK_2_470(net730_c1,net730);
INTERCONNECT SplitCLK_4_288_SplitCLK_4_287(net731_c1,net731);
INTERCONNECT SplitCLK_4_287_AND2T_84_n108(net732_c1,net732);
INTERCONNECT SplitCLK_4_287_DFFT_175__FPB_n565(net733_c1,net733);
INTERCONNECT SplitCLK_6_286_SplitCLK_4_284(net734_c1,net734);
INTERCONNECT SplitCLK_6_286_SplitCLK_4_285(net735_c1,net735);
INTERCONNECT SplitCLK_4_285_AND2T_76_n100(net736_c1,net736);
INTERCONNECT SplitCLK_4_285_OR2T_79_n103(net737_c1,net737);
INTERCONNECT SplitCLK_4_284_OR2T_72_n96(net738_c1,net738);
INTERCONNECT SplitCLK_4_284_DFFT_191__FPB_n581(net739_c1,net739);
INTERCONNECT SplitCLK_4_283_SplitCLK_4_280(net740_c1,net740);
INTERCONNECT SplitCLK_4_283_SplitCLK_2_282(net741_c1,net741);
INTERCONNECT SplitCLK_2_282_SplitCLK_2_456(net742_c1,net742);
INTERCONNECT SplitCLK_2_282_SplitCLK_4_281(net743_c1,net743);
INTERCONNECT SplitCLK_4_281_OR2T_90_n114(net744_c1,net744);
INTERCONNECT SplitCLK_4_281_DFFT_193__FPB_n583(net745_c1,net745);
INTERCONNECT SplitCLK_4_280_SplitCLK_4_278(net746_c1,net746);
INTERCONNECT SplitCLK_4_280_SplitCLK_4_279(net747_c1,net747);
INTERCONNECT SplitCLK_4_279_OR2T_73_n97(net748_c1,net748);
INTERCONNECT SplitCLK_4_279_OR2T_88_n112(net749_c1,net749);
INTERCONNECT SplitCLK_4_278_OR2T_89_n113(net750_c1,net750);
INTERCONNECT SplitCLK_4_278_DFFT_178__FPB_n568(net751_c1,net751);
INTERCONNECT SplitCLK_6_277_SplitCLK_0_249(net752_c1,net752);
INTERCONNECT SplitCLK_6_277_SplitCLK_2_276(net753_c1,net753);
INTERCONNECT SplitCLK_2_276_SplitCLK_6_262(net754_c1,net754);
INTERCONNECT SplitCLK_2_276_SplitCLK_4_275(net755_c1,net755);
INTERCONNECT SplitCLK_4_275_SplitCLK_0_268(net756_c1,net756);
INTERCONNECT SplitCLK_4_275_SplitCLK_2_274(net757_c1,net757);
INTERCONNECT SplitCLK_2_274_SplitCLK_6_271(net758_c1,net758);
INTERCONNECT SplitCLK_2_274_SplitCLK_4_273(net759_c1,net759);
INTERCONNECT SplitCLK_4_273_SplitCLK_2_450(net760_c1,net760);
INTERCONNECT SplitCLK_4_273_SplitCLK_4_272(net761_c1,net761);
INTERCONNECT SplitCLK_4_272_AND2T_41_n65(net762_c1,net762);
INTERCONNECT SplitCLK_4_272_AND2T_44_n68(net763_c1,net763);
INTERCONNECT SplitCLK_6_271_SplitCLK_4_269(net764_c1,net764);
INTERCONNECT SplitCLK_6_271_SplitCLK_4_270(net765_c1,net765);
INTERCONNECT SplitCLK_4_270_AND2T_20_n44(net766_c1,net766);
INTERCONNECT SplitCLK_4_270_OR2T_16_n40(net767_c1,net767);
INTERCONNECT SplitCLK_4_269_OR2T_27_n51(net768_c1,net768);
INTERCONNECT SplitCLK_4_269_DFFT_120__FPB_n510(net769_c1,net769);
INTERCONNECT SplitCLK_0_268_SplitCLK_6_265(net770_c1,net770);
INTERCONNECT SplitCLK_0_268_SplitCLK_4_267(net771_c1,net771);
INTERCONNECT SplitCLK_4_267_SplitCLK_2_444(net772_c1,net772);
INTERCONNECT SplitCLK_4_267_SplitCLK_4_266(net773_c1,net773);
INTERCONNECT SplitCLK_4_266_AND2T_61_n85(net774_c1,net774);
INTERCONNECT SplitCLK_4_266_AND2T_58_n82(net775_c1,net775);
INTERCONNECT SplitCLK_6_265_SplitCLK_4_263(net776_c1,net776);
INTERCONNECT SplitCLK_6_265_SplitCLK_4_264(net777_c1,net777);
INTERCONNECT SplitCLK_4_264_AND2T_26_n50(net778_c1,net778);
INTERCONNECT SplitCLK_4_264_DFFT_126__FPB_n516(net779_c1,net779);
INTERCONNECT SplitCLK_4_263_AND2T_30_n54(net780_c1,net780);
INTERCONNECT SplitCLK_4_263_OR2T_33_n57(net781_c1,net781);
INTERCONNECT SplitCLK_6_262_SplitCLK_6_255(net782_c1,net782);
INTERCONNECT SplitCLK_6_262_SplitCLK_6_261(net783_c1,net783);
INTERCONNECT SplitCLK_6_261_SplitCLK_6_258(net784_c1,net784);
INTERCONNECT SplitCLK_6_261_SplitCLK_4_260(net785_c1,net785);
INTERCONNECT SplitCLK_4_260_SplitCLK_2_455(net786_c1,net786);
INTERCONNECT SplitCLK_4_260_SplitCLK_4_259(net787_c1,net787);
INTERCONNECT SplitCLK_4_259_AND2T_22_n46(net788_c1,net788);
INTERCONNECT SplitCLK_4_259_AND2T_24_n48(net789_c1,net789);
INTERCONNECT SplitCLK_6_258_SplitCLK_4_256(net790_c1,net790);
INTERCONNECT SplitCLK_6_258_SplitCLK_4_257(net791_c1,net791);
INTERCONNECT SplitCLK_4_257_DFFT_222__FPB_n612(net792_c1,net792);
INTERCONNECT SplitCLK_4_257_NOTT_97_n130(net793_c1,net793);
INTERCONNECT SplitCLK_4_256_AND2T_14_n38(net794_c1,net794);
INTERCONNECT SplitCLK_4_256_DFFT_221__FPB_n611(net795_c1,net795);
INTERCONNECT SplitCLK_6_255_SplitCLK_6_252(net796_c1,net796);
INTERCONNECT SplitCLK_6_255_SplitCLK_0_254(net797_c1,net797);
INTERCONNECT SplitCLK_0_254_SplitCLK_2_454(net798_c1,net798);
INTERCONNECT SplitCLK_0_254_SplitCLK_4_253(net799_c1,net799);
INTERCONNECT SplitCLK_4_253_AND2T_15_n39(net800_c1,net800);
INTERCONNECT SplitCLK_4_253_DFFT_117__FPB_n507(net801_c1,net801);
INTERCONNECT SplitCLK_6_252_SplitCLK_4_250(net802_c1,net802);
INTERCONNECT SplitCLK_6_252_SplitCLK_4_251(net803_c1,net803);
INTERCONNECT SplitCLK_4_251_DFFT_220__FPB_n610(net804_c1,net804);
INTERCONNECT SplitCLK_4_251_DFFT_219__FPB_n609(net805_c1,net805);
INTERCONNECT SplitCLK_4_250_DFFT_229_state_obs3(net806_c1,net806);
INTERCONNECT SplitCLK_4_250_DFFT_102__PIPL_n138(net807_c1,net807);
INTERCONNECT SplitCLK_0_249_SplitCLK_6_235(net808_c1,net808);
INTERCONNECT SplitCLK_0_249_SplitCLK_4_248(net809_c1,net809);
INTERCONNECT SplitCLK_4_248_SplitCLK_4_241(net810_c1,net810);
INTERCONNECT SplitCLK_4_248_SplitCLK_2_247(net811_c1,net811);
INTERCONNECT SplitCLK_2_247_SplitCLK_6_244(net812_c1,net812);
INTERCONNECT SplitCLK_2_247_SplitCLK_2_246(net813_c1,net813);
INTERCONNECT SplitCLK_2_246_SplitCLK_2_452(net814_c1,net814);
INTERCONNECT SplitCLK_2_246_SplitCLK_4_245(net815_c1,net815);
INTERCONNECT SplitCLK_4_245_AND2T_74_n98(net816_c1,net816);
INTERCONNECT SplitCLK_4_245_OR2T_59_n83(net817_c1,net817);
INTERCONNECT SplitCLK_6_244_SplitCLK_0_242(net818_c1,net818);
INTERCONNECT SplitCLK_6_244_SplitCLK_4_243(net819_c1,net819);
INTERCONNECT SplitCLK_4_243_DFFT_161__FPB_n551(net820_c1,net820);
INTERCONNECT SplitCLK_4_243_DFFT_173__FPB_n563(net821_c1,net821);
INTERCONNECT SplitCLK_0_242_AND2T_32_n56(net822_c1,net822);
INTERCONNECT SplitCLK_0_242_DFFT_176__FPB_n566(net823_c1,net823);
INTERCONNECT SplitCLK_4_241_SplitCLK_6_238(net824_c1,net824);
INTERCONNECT SplitCLK_4_241_SplitCLK_4_240(net825_c1,net825);
INTERCONNECT SplitCLK_4_240_SplitCLK_2_449(net826_c1,net826);
INTERCONNECT SplitCLK_4_240_SplitCLK_4_239(net827_c1,net827);
INTERCONNECT SplitCLK_4_239_AND2T_62_n86(net828_c1,net828);
INTERCONNECT SplitCLK_4_239_DFFT_160__FPB_n550(net829_c1,net829);
INTERCONNECT SplitCLK_6_238_SplitCLK_4_236(net830_c1,net830);
INTERCONNECT SplitCLK_6_238_SplitCLK_4_237(net831_c1,net831);
INTERCONNECT SplitCLK_4_237_AND2T_86_n110(net832_c1,net832);
INTERCONNECT SplitCLK_4_237_DFFT_192__FPB_n582(net833_c1,net833);
INTERCONNECT SplitCLK_4_236_AND2T_63_n87(net834_c1,net834);
INTERCONNECT SplitCLK_4_236_DFFT_127__FPB_n517(net835_c1,net835);
INTERCONNECT SplitCLK_6_235_SplitCLK_0_228(net836_c1,net836);
INTERCONNECT SplitCLK_6_235_SplitCLK_6_234(net837_c1,net837);
INTERCONNECT SplitCLK_6_234_SplitCLK_6_231(net838_c1,net838);
INTERCONNECT SplitCLK_6_234_SplitCLK_4_233(net839_c1,net839);
INTERCONNECT SplitCLK_4_233_SplitCLK_2_467(net840_c1,net840);
INTERCONNECT SplitCLK_4_233_SplitCLK_4_232(net841_c1,net841);
INTERCONNECT SplitCLK_4_232_AND2T_77_n101(net842_c1,net842);
INTERCONNECT SplitCLK_4_232_DFFT_140__FPB_n530(net843_c1,net843);
INTERCONNECT SplitCLK_6_231_SplitCLK_4_229(net844_c1,net844);
INTERCONNECT SplitCLK_6_231_SplitCLK_4_230(net845_c1,net845);
INTERCONNECT SplitCLK_4_230_DFFT_218__FPB_n608(net846_c1,net846);
INTERCONNECT SplitCLK_4_230_DFFT_228__FPB_n618(net847_c1,net847);
INTERCONNECT SplitCLK_4_229_DFFT_103__PIPL_n139(net848_c1,net848);
INTERCONNECT SplitCLK_4_229_DFFT_227__FPB_n617(net849_c1,net849);
INTERCONNECT SplitCLK_0_228_SplitCLK_6_225(net850_c1,net850);
INTERCONNECT SplitCLK_0_228_SplitCLK_2_227(net851_c1,net851);
INTERCONNECT SplitCLK_2_227_SplitCLK_2_460(net852_c1,net852);
INTERCONNECT SplitCLK_2_227_SplitCLK_4_226(net853_c1,net853);
INTERCONNECT SplitCLK_4_226_DFFT_110__FBL_n500(net854_c1,net854);
INTERCONNECT SplitCLK_4_226_DFFT_113__FPB_n503(net855_c1,net855);
INTERCONNECT SplitCLK_6_225_SplitCLK_4_223(net856_c1,net856);
INTERCONNECT SplitCLK_6_225_SplitCLK_4_224(net857_c1,net857);
INTERCONNECT SplitCLK_4_224_DFFT_224__FPB_n614(net858_c1,net858);
INTERCONNECT SplitCLK_4_224_DFFT_225__FPB_n615(net859_c1,net859);
INTERCONNECT SplitCLK_4_223_DFFT_115__FPB_n505(net860_c1,net860);
INTERCONNECT SplitCLK_4_223_DFFT_226__FPB_n616(net861_c1,net861);
INTERCONNECT GCLK_Pad_SplitCLK_0_477(GCLK_Pad,net862);
INTERCONNECT Split_HOLD_566_DFFT_137__FPB_n527(net863_c1,net863);
INTERCONNECT Split_HOLD_567_DFFT_214__FPB_n604(net864_c1,net864);
INTERCONNECT Split_HOLD_568_NOTT_97_n130(net865_c1,net865);
INTERCONNECT Split_HOLD_569_DFFT_125__FPB_n515(net866_c1,net866);
INTERCONNECT Split_HOLD_570_DFFT_204__FPB_n594(net867_c1,net867);
INTERCONNECT Split_HOLD_571_DFFT_123__FPB_n513(net868_c1,net868);

endmodule
