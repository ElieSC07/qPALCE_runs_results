module TAP_route(
input GCLK_Pad,
input TMS_Pad,
input TRST_Pad,
output state_obs0_Pad,
output state_obs1_Pad,
output state_obs2_Pad,
output state_obs3_Pad);

wire TMS_Pad;
wire net0;
wire net1_c1;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire TRST_Pad;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire net266;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire state_obs0_Pad;
wire net437_c1;
wire state_obs1_Pad;
wire net438_c1;
wire state_obs2_Pad;
wire net439_c1;
wire state_obs3_Pad;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire net486_c1;
wire net486;
wire net487_c1;
wire net487;
wire net488_c1;
wire net488;
wire net489_c1;
wire net489;
wire net490_c1;
wire net490;
wire net491_c1;
wire net491;
wire net492_c1;
wire net492;
wire net493_c1;
wire net493;
wire net494_c1;
wire net494;
wire net495_c1;
wire net495;
wire net496_c1;
wire net496;
wire net497_c1;
wire net497;
wire net498_c1;
wire net498;
wire net499_c1;
wire net499;
wire net500_c1;
wire net500;
wire net501_c1;
wire net501;
wire net502_c1;
wire net502;
wire net503_c1;
wire net503;
wire net504_c1;
wire net504;
wire net505_c1;
wire net505;
wire net506_c1;
wire net506;
wire net507_c1;
wire net507;
wire net508_c1;
wire net508;
wire net509_c1;
wire net509;
wire net510_c1;
wire net510;
wire net511_c1;
wire net511;
wire net512_c1;
wire net512;
wire net513_c1;
wire net513;
wire net514_c1;
wire net514;
wire net515_c1;
wire net515;
wire net516_c1;
wire net516;
wire net517_c1;
wire net517;
wire net518_c1;
wire net518;
wire net519_c1;
wire net519;
wire net520_c1;
wire net520;
wire net521_c1;
wire net521;
wire net522_c1;
wire net522;
wire net523_c1;
wire net523;
wire net524_c1;
wire net524;
wire net525_c1;
wire net525;
wire net526_c1;
wire net526;
wire net527_c1;
wire net527;
wire net528_c1;
wire net528;
wire net529_c1;
wire net529;
wire net530_c1;
wire net530;
wire net531_c1;
wire net531;
wire net532_c1;
wire net532;
wire net533_c1;
wire net533;
wire net534_c1;
wire net534;
wire net535_c1;
wire net535;
wire net536_c1;
wire net536;
wire net537_c1;
wire net537;
wire net538_c1;
wire net538;
wire net539_c1;
wire net539;
wire net540_c1;
wire net540;
wire net541_c1;
wire net541;
wire net542_c1;
wire net542;
wire net543_c1;
wire net543;
wire net544_c1;
wire net544;
wire net545_c1;
wire net545;
wire net546_c1;
wire net546;
wire net547_c1;
wire net547;
wire net548_c1;
wire net548;
wire net549_c1;
wire net549;
wire net550_c1;
wire net550;
wire net551_c1;
wire net551;
wire net552_c1;
wire net552;
wire net553_c1;
wire net553;
wire net554_c1;
wire net554;
wire net555_c1;
wire net555;
wire net556_c1;
wire net556;
wire net557_c1;
wire net557;
wire net558_c1;
wire net558;
wire net559_c1;
wire net559;
wire net560_c1;
wire net560;
wire net561_c1;
wire net561;
wire net562_c1;
wire net562;
wire net563_c1;
wire net563;
wire net564_c1;
wire net564;
wire net565_c1;
wire net565;
wire net566_c1;
wire net566;
wire net567_c1;
wire net567;
wire net568_c1;
wire net568;
wire net569_c1;
wire net569;
wire net570_c1;
wire net570;
wire net571_c1;
wire net571;
wire net572_c1;
wire net572;
wire net573_c1;
wire net573;
wire net574_c1;
wire net574;
wire net575_c1;
wire net575;
wire net576_c1;
wire net576;
wire net577_c1;
wire net577;
wire net578_c1;
wire net578;
wire net579_c1;
wire net579;
wire net580_c1;
wire net580;
wire net581_c1;
wire net581;
wire net582_c1;
wire net582;
wire net583_c1;
wire net583;
wire net584_c1;
wire net584;
wire net585_c1;
wire net585;
wire net586_c1;
wire net586;
wire net587_c1;
wire net587;
wire net588_c1;
wire net588;
wire net589_c1;
wire net589;
wire net590_c1;
wire net590;
wire net591_c1;
wire net591;
wire net592_c1;
wire net592;
wire net593_c1;
wire net593;
wire net594_c1;
wire net594;
wire net595_c1;
wire net595;
wire net596_c1;
wire net596;
wire net597_c1;
wire net597;
wire net598_c1;
wire net598;
wire net599_c1;
wire net599;
wire net600_c1;
wire net600;
wire net601_c1;
wire net601;
wire net602_c1;
wire net602;
wire net603_c1;
wire net603;
wire net604_c1;
wire net604;
wire net605_c1;
wire net605;
wire net606_c1;
wire net606;
wire net607_c1;
wire net607;
wire net608_c1;
wire net608;
wire net609_c1;
wire net609;
wire net610_c1;
wire net610;
wire net611_c1;
wire net611;
wire net612_c1;
wire net612;
wire net613_c1;
wire net613;
wire net614_c1;
wire net614;
wire net615_c1;
wire net615;
wire net616_c1;
wire net616;
wire net617_c1;
wire net617;
wire net618_c1;
wire net618;
wire net619_c1;
wire net619;
wire net620_c1;
wire net620;
wire net621_c1;
wire net621;
wire net622_c1;
wire net622;
wire net623_c1;
wire net623;
wire net624_c1;
wire net624;
wire net625_c1;
wire net625;
wire net626_c1;
wire net626;
wire net627_c1;
wire net627;
wire net628_c1;
wire net628;
wire net629_c1;
wire net629;
wire net630_c1;
wire net630;
wire net631_c1;
wire net631;
wire net632_c1;
wire net632;
wire net633_c1;
wire net633;
wire net634_c1;
wire net634;
wire net635_c1;
wire net635;
wire net636_c1;
wire net636;
wire net637_c1;
wire net637;
wire net638_c1;
wire net638;
wire net639_c1;
wire net639;
wire net640_c1;
wire net640;
wire net641_c1;
wire net641;
wire net642_c1;
wire net642;
wire net643_c1;
wire net643;
wire net644_c1;
wire net644;
wire net645_c1;
wire net645;
wire net646_c1;
wire net646;
wire net647_c1;
wire net647;
wire net648_c1;
wire net648;
wire net649_c1;
wire net649;
wire net650_c1;
wire net650;
wire net651_c1;
wire net651;
wire net652_c1;
wire net652;
wire net653_c1;
wire net653;
wire net654_c1;
wire net654;
wire net655_c1;
wire net655;
wire net656_c1;
wire net656;
wire net657_c1;
wire net657;
wire net658_c1;
wire net658;
wire net659_c1;
wire net659;
wire net660_c1;
wire net660;
wire net661_c1;
wire net661;
wire net662_c1;
wire net662;
wire net663_c1;
wire net663;
wire net664_c1;
wire net664;
wire net665_c1;
wire net665;
wire net666_c1;
wire net666;
wire net667_c1;
wire net667;
wire net668_c1;
wire net668;
wire net669_c1;
wire net669;
wire net670_c1;
wire net670;
wire net671_c1;
wire net671;
wire net672_c1;
wire net672;
wire net673_c1;
wire net673;
wire net674_c1;
wire net674;
wire net675_c1;
wire net675;
wire net676_c1;
wire net676;
wire net677_c1;
wire net677;
wire net678_c1;
wire net678;
wire net679_c1;
wire net679;
wire net680_c1;
wire net680;
wire net681_c1;
wire net681;
wire net682_c1;
wire net682;
wire net683_c1;
wire net683;
wire net684_c1;
wire net684;
wire net685_c1;
wire net685;
wire net686_c1;
wire net686;
wire net687_c1;
wire net687;
wire net688_c1;
wire net688;
wire net689_c1;
wire net689;
wire net690_c1;
wire net690;
wire net691_c1;
wire net691;
wire net692_c1;
wire net692;
wire net693_c1;
wire net693;
wire net694_c1;
wire net694;
wire net695_c1;
wire net695;
wire net696_c1;
wire net696;
wire net697_c1;
wire net697;
wire net698_c1;
wire net698;
wire net699_c1;
wire net699;
wire net700_c1;
wire net700;
wire net701_c1;
wire net701;
wire net702_c1;
wire net702;
wire net703_c1;
wire net703;
wire net704_c1;
wire net704;
wire net705_c1;
wire net705;
wire net706_c1;
wire net706;
wire net707_c1;
wire net707;
wire net708_c1;
wire net708;
wire net709_c1;
wire net709;
wire net710_c1;
wire net710;
wire net711_c1;
wire net711;
wire net712_c1;
wire net712;
wire net713_c1;
wire net713;
wire net714_c1;
wire net714;
wire net715_c1;
wire net715;
wire net716_c1;
wire net716;
wire net717_c1;
wire net717;
wire net718_c1;
wire net718;
wire net719_c1;
wire net719;
wire net720_c1;
wire net720;
wire net721_c1;
wire net721;
wire net722_c1;
wire net722;
wire net723_c1;
wire net723;
wire net724_c1;
wire net724;
wire net725_c1;
wire net725;
wire net726_c1;
wire net726;
wire net727_c1;
wire net727;
wire net728_c1;
wire net728;
wire net729_c1;
wire net729;
wire net730_c1;
wire net730;
wire net731_c1;
wire net731;
wire net732_c1;
wire net732;
wire net733_c1;
wire net733;
wire net734_c1;
wire net734;
wire net735_c1;
wire net735;
wire net736_c1;
wire net736;
wire net737_c1;
wire net737;
wire net738_c1;
wire net738;
wire net739_c1;
wire net739;
wire net740_c1;
wire net740;
wire net741_c1;
wire net741;
wire net742_c1;
wire net742;
wire net743_c1;
wire net743;
wire net744_c1;
wire net744;
wire net745_c1;
wire net745;
wire net746_c1;
wire net746;
wire net747_c1;
wire net747;
wire net748_c1;
wire net748;
wire net749_c1;
wire net749;
wire net750_c1;
wire net750;
wire net751_c1;
wire net751;
wire net752_c1;
wire net752;
wire net753_c1;
wire net753;
wire net754_c1;
wire net754;
wire net755_c1;
wire net755;
wire net756_c1;
wire net756;
wire net757_c1;
wire net757;
wire net758_c1;
wire net758;
wire net759_c1;
wire net759;
wire net760_c1;
wire net760;
wire net761_c1;
wire net761;
wire net762_c1;
wire net762;
wire net763_c1;
wire net763;
wire net764_c1;
wire net764;
wire net765_c1;
wire net765;
wire net766_c1;
wire net766;
wire net767_c1;
wire net767;
wire net768_c1;
wire net768;
wire net769_c1;
wire net769;
wire net770_c1;
wire net770;
wire net771_c1;
wire net771;
wire net772_c1;
wire net772;
wire net773_c1;
wire net773;
wire net774_c1;
wire net774;
wire net775_c1;
wire net775;
wire net776_c1;
wire net776;
wire net777_c1;
wire net777;
wire net778_c1;
wire net778;
wire net779_c1;
wire net779;
wire net780_c1;
wire net780;
wire net781_c1;
wire net781;
wire net782_c1;
wire net782;
wire net783_c1;
wire net783;
wire net784_c1;
wire net784;
wire net785_c1;
wire net785;
wire net786_c1;
wire net786;
wire net787_c1;
wire net787;
wire net788_c1;
wire net788;
wire net789_c1;
wire net789;
wire net790_c1;
wire net790;
wire net791_c1;
wire net791;
wire net792_c1;
wire net792;
wire net793_c1;
wire net793;
wire net794_c1;
wire net794;
wire net795_c1;
wire net795;
wire net796_c1;
wire net796;
wire net797_c1;
wire net797;
wire net798_c1;
wire net798;
wire net799_c1;
wire net799;
wire net800_c1;
wire net800;
wire net801_c1;
wire net801;
wire net802_c1;
wire net802;
wire net803_c1;
wire net803;
wire net804_c1;
wire net804;
wire net805_c1;
wire net805;
wire net806_c1;
wire net806;
wire net807_c1;
wire net807;
wire net808_c1;
wire net808;
wire net809_c1;
wire net809;
wire net810_c1;
wire net810;
wire net811_c1;
wire net811;
wire net812_c1;
wire net812;
wire net813_c1;
wire net813;
wire net814_c1;
wire net814;
wire net815_c1;
wire net815;
wire net816_c1;
wire net816;
wire net817_c1;
wire net817;
wire net818_c1;
wire net818;
wire net819_c1;
wire net819;
wire net820_c1;
wire net820;
wire net821_c1;
wire net821;
wire net822_c1;
wire net822;
wire net823_c1;
wire net823;
wire net824_c1;
wire net824;
wire net825_c1;
wire net825;
wire net826_c1;
wire net826;
wire net827_c1;
wire net827;
wire net828_c1;
wire net828;
wire net829_c1;
wire net829;
wire net830_c1;
wire net830;
wire net831_c1;
wire net831;
wire net832_c1;
wire net832;
wire net833_c1;
wire net833;
wire net834_c1;
wire net834;
wire net835_c1;
wire net835;
wire net836_c1;
wire net836;
wire net837_c1;
wire net837;
wire net838_c1;
wire net838;
wire net839_c1;
wire net839;
wire net840_c1;
wire net840;
wire net841_c1;
wire net841;
wire net842_c1;
wire net842;
wire net843_c1;
wire net843;
wire net844_c1;
wire net844;
wire net845_c1;
wire net845;
wire net846_c1;
wire net846;
wire net847_c1;
wire net847;
wire net848_c1;
wire net848;
wire net849_c1;
wire net849;
wire net850_c1;
wire net850;
wire net851_c1;
wire net851;
wire net852_c1;
wire net852;
wire net853_c1;
wire net853;
wire net854_c1;
wire net854;
wire net855_c1;
wire net855;
wire net856_c1;
wire net856;
wire net857_c1;
wire net857;
wire net858_c1;
wire net858;
wire net859_c1;
wire net859;
wire net860_c1;
wire net860;
wire net861_c1;
wire net861;
wire net862_c1;
wire net862;
wire net863_c1;
wire net863;
wire net864_c1;
wire net864;
wire net865_c1;
wire net865;
wire net866_c1;
wire net866;
wire net867_c1;
wire net867;
wire net868_c1;
wire net868;
wire net869_c1;
wire net869;
wire net870_c1;
wire net870;
wire net871_c1;
wire net871;
wire net872_c1;
wire net872;
wire net873_c1;
wire net873;
wire net874_c1;
wire net874;
wire net875_c1;
wire net875;
wire net876_c1;
wire net876;
wire net877_c1;
wire net877;
wire net878_c1;
wire net878;
wire net879_c1;
wire net879;
wire net880_c1;
wire net880;
wire net881_c1;
wire net881;
wire net882_c1;
wire net882;
wire net883_c1;
wire net883;
wire net884_c1;
wire net884;
wire net885_c1;
wire net885;
wire net886_c1;
wire net886;
wire net887_c1;
wire net887;
wire net888_c1;
wire net888;
wire net889_c1;
wire net889;
wire net890_c1;
wire net890;
wire net891_c1;
wire net891;
wire net892_c1;
wire net892;
wire net893_c1;
wire net893;
wire net894_c1;
wire net894;
wire net895_c1;
wire net895;
wire net896_c1;
wire net896;
wire net897_c1;
wire net897;
wire net898_c1;
wire net898;
wire net899_c1;
wire net899;
wire net900_c1;
wire net900;
wire net901_c1;
wire net901;
wire net902_c1;
wire net902;
wire net903_c1;
wire net903;
wire net904_c1;
wire net904;
wire net905_c1;
wire net905;
wire net906_c1;
wire net906;
wire net907_c1;
wire net907;
wire net908_c1;
wire net908;
wire net909_c1;
wire net909;
wire net910_c1;
wire net910;
wire net911_c1;
wire net911;
wire net912_c1;
wire net912;
wire net913_c1;
wire net913;
wire net914_c1;
wire net914;
wire net915_c1;
wire net915;
wire net916_c1;
wire net916;
wire net917_c1;
wire net917;
wire net918_c1;
wire net918;
wire net919_c1;
wire net919;
wire net920_c1;
wire net920;
wire net921_c1;
wire net921;
wire net922_c1;
wire net922;
wire net923_c1;
wire net923;
wire net924_c1;
wire net924;
wire net925_c1;
wire net925;
wire net926_c1;
wire net926;
wire net927_c1;
wire net927;
wire net928_c1;
wire net928;
wire net929_c1;
wire net929;
wire net930_c1;
wire net930;
wire net931_c1;
wire net931;
wire net932_c1;
wire net932;
wire net933_c1;
wire net933;
wire net934_c1;
wire net934;
wire net935_c1;
wire net935;
wire net936_c1;
wire net936;
wire net937_c1;
wire net937;
wire net938_c1;
wire net938;
wire net939_c1;
wire net939;
wire net940_c1;
wire net940;
wire net941_c1;
wire net941;
wire net942_c1;
wire net942;
wire net943_c1;
wire net943;
wire net944_c1;
wire net944;
wire net945_c1;
wire net945;
wire net946_c1;
wire net946;
wire net947_c1;
wire net947;
wire net948_c1;
wire net948;
wire net949_c1;
wire net949;
wire net950_c1;
wire net950;
wire net951_c1;
wire net951;
wire net952_c1;
wire net952;
wire net953_c1;
wire net953;
wire net954_c1;
wire net954;
wire net955_c1;
wire net955;
wire net956_c1;
wire net956;
wire net957_c1;
wire net957;
wire net958_c1;
wire net958;
wire net959_c1;
wire net959;
wire net960_c1;
wire net960;
wire net961_c1;
wire net961;
wire net962_c1;
wire net962;
wire net963_c1;
wire net963;
wire net964_c1;
wire net964;
wire net965_c1;
wire net965;
wire net966_c1;
wire net966;
wire net967_c1;
wire net967;
wire net968_c1;
wire net968;
wire net969_c1;
wire net969;
wire net970_c1;
wire net970;
wire net971_c1;
wire net971;
wire net972_c1;
wire net972;
wire net973_c1;
wire net973;
wire net974_c1;
wire net974;
wire net975_c1;
wire net975;
wire net976_c1;
wire net976;
wire net977_c1;
wire net977;
wire net978_c1;
wire net978;
wire net979_c1;
wire net979;
wire net980_c1;
wire net980;
wire net981_c1;
wire net981;
wire net982_c1;
wire net982;
wire net983_c1;
wire net983;
wire net984_c1;
wire net984;
wire net985_c1;
wire net985;
wire net986_c1;
wire net986;
wire net987_c1;
wire net987;
wire net988_c1;
wire net988;
wire net989_c1;
wire net989;
wire net990_c1;
wire net990;
wire net991_c1;
wire net991;
wire net992_c1;
wire net992;
wire net993_c1;
wire net993;
wire net994_c1;
wire net994;
wire net995_c1;
wire net995;
wire net996_c1;
wire net996;
wire net997_c1;
wire net997;
wire net998_c1;
wire net998;
wire net999_c1;
wire net999;
wire net1000_c1;
wire net1000;
wire net1001_c1;
wire net1001;
wire net1002_c1;
wire net1002;
wire net1003_c1;
wire net1003;
wire net1004_c1;
wire net1004;
wire net1005_c1;
wire net1005;
wire net1006_c1;
wire net1006;
wire net1007_c1;
wire net1007;
wire net1008_c1;
wire net1008;
wire net1009_c1;
wire net1009;
wire net1010_c1;
wire net1010;
wire net1011_c1;
wire net1011;
wire net1012_c1;
wire net1012;
wire net1013_c1;
wire net1013;
wire net1014_c1;
wire net1014;
wire net1015_c1;
wire net1015;
wire net1016_c1;
wire net1016;
wire net1017_c1;
wire net1017;
wire net1018_c1;
wire net1018;
wire net1019_c1;
wire net1019;
wire net1020_c1;
wire net1020;
wire net1021_c1;
wire net1021;
wire net1022_c1;
wire net1022;
wire net1023_c1;
wire net1023;
wire net1024_c1;
wire net1024;
wire net1025_c1;
wire net1025;
wire net1026_c1;
wire net1026;
wire net1027_c1;
wire net1027;
wire net1028_c1;
wire net1028;
wire net1029_c1;
wire net1029;
wire net1030_c1;
wire net1030;
wire net1031_c1;
wire net1031;
wire net1032_c1;
wire net1032;
wire net1033_c1;
wire net1033;
wire net1034_c1;
wire net1034;
wire net1035_c1;
wire net1035;
wire net1036_c1;
wire net1036;
wire net1037_c1;
wire net1037;
wire net1038_c1;
wire net1038;
wire net1039_c1;
wire net1039;
wire net1040_c1;
wire net1040;
wire net1041_c1;
wire net1041;
wire net1042_c1;
wire net1042;
wire net1043_c1;
wire net1043;
wire net1044_c1;
wire net1044;
wire net1045_c1;
wire net1045;
wire net1046_c1;
wire net1046;
wire net1047_c1;
wire net1047;
wire net1048_c1;
wire net1048;
wire net1049_c1;
wire net1049;
wire net1050_c1;
wire net1050;
wire net1051_c1;
wire net1051;
wire net1052_c1;
wire net1052;
wire net1053_c1;
wire net1053;
wire net1054_c1;
wire net1054;
wire net1055_c1;
wire net1055;
wire net1056_c1;
wire net1056;
wire net1057_c1;
wire net1057;
wire net1058_c1;
wire net1058;
wire net1059_c1;
wire net1059;
wire net1060_c1;
wire net1060;
wire net1061_c1;
wire net1061;
wire net1062_c1;
wire net1062;
wire net1063_c1;
wire net1063;
wire net1064_c1;
wire net1064;
wire net1065_c1;
wire net1065;
wire net1066_c1;
wire net1066;
wire net1067_c1;
wire net1067;
wire net1068_c1;
wire net1068;
wire net1069_c1;
wire net1069;
wire net1070_c1;
wire net1070;
wire net1071_c1;
wire net1071;
wire net1072_c1;
wire net1072;
wire net1073_c1;
wire net1073;
wire net1074_c1;
wire net1074;
wire net1075_c1;
wire net1075;
wire net1076_c1;
wire net1076;
wire net1077_c1;
wire net1077;
wire net1078_c1;
wire net1078;
wire net1079_c1;
wire net1079;
wire net1080_c1;
wire net1080;
wire net1081_c1;
wire net1081;
wire net1082_c1;
wire net1082;
wire net1083_c1;
wire net1083;
wire net1084_c1;
wire net1084;
wire net1085_c1;
wire net1085;
wire net1086_c1;
wire net1086;
wire net1087_c1;
wire net1087;
wire net1088_c1;
wire net1088;
wire net1089_c1;
wire net1089;
wire net1090_c1;
wire net1090;
wire net1091_c1;
wire net1091;
wire net1092_c1;
wire net1092;
wire net1093_c1;
wire net1093;
wire net1094_c1;
wire net1094;
wire net1095_c1;
wire net1095;
wire net1096_c1;
wire net1096;
wire net1097_c1;
wire net1097;
wire net1098_c1;
wire net1098;
wire net1099_c1;
wire net1099;
wire net1100_c1;
wire net1100;
wire net1101_c1;
wire net1101;
wire net1102_c1;
wire net1102;
wire net1103_c1;
wire net1103;
wire net1104_c1;
wire net1104;
wire net1105_c1;
wire net1105;
wire net1106_c1;
wire net1106;
wire net1107_c1;
wire net1107;
wire net1108_c1;
wire net1108;
wire net1109_c1;
wire net1109;
wire net1110_c1;
wire net1110;
wire net1111_c1;
wire net1111;
wire net1112_c1;
wire net1112;
wire net1113_c1;
wire net1113;
wire net1114_c1;
wire net1114;
wire net1115_c1;
wire net1115;
wire net1116_c1;
wire net1116;
wire net1117_c1;
wire net1117;
wire net1118_c1;
wire net1118;
wire net1119_c1;
wire net1119;
wire net1120_c1;
wire net1120;
wire net1121_c1;
wire net1121;
wire net1122_c1;
wire net1122;
wire net1123_c1;
wire net1123;
wire net1124_c1;
wire net1124;
wire net1125_c1;
wire net1125;
wire net1126_c1;
wire net1126;
wire net1127_c1;
wire net1127;
wire net1128_c1;
wire net1128;
wire net1129_c1;
wire net1129;
wire net1130_c1;
wire net1130;
wire net1131_c1;
wire net1131;
wire net1132_c1;
wire net1132;
wire net1133_c1;
wire net1133;
wire net1134_c1;
wire net1134;
wire net1135_c1;
wire net1135;
wire net1136_c1;
wire net1136;
wire net1137_c1;
wire net1137;
wire net1138_c1;
wire net1138;
wire net1139_c1;
wire net1139;
wire net1140_c1;
wire net1140;
wire net1141_c1;
wire net1141;
wire net1142_c1;
wire net1142;
wire net1143_c1;
wire net1143;
wire net1144_c1;
wire net1144;
wire net1145_c1;
wire net1145;
wire net1146_c1;
wire net1146;
wire net1147_c1;
wire net1147;
wire net1148_c1;
wire net1148;
wire net1149_c1;
wire net1149;
wire net1150_c1;
wire net1150;
wire net1151_c1;
wire net1151;
wire net1152_c1;
wire net1152;
wire net1153_c1;
wire net1153;
wire net1154_c1;
wire net1154;
wire net1155_c1;
wire net1155;
wire net1156_c1;
wire net1156;
wire net1157_c1;
wire net1157;
wire net1158_c1;
wire net1158;
wire net1159_c1;
wire net1159;
wire net1160_c1;
wire net1160;
wire net1161_c1;
wire net1161;
wire net1162_c1;
wire net1162;
wire net1163_c1;
wire net1163;
wire net1164_c1;
wire net1164;
wire net1165_c1;
wire net1165;
wire net1166_c1;
wire net1166;
wire net1167_c1;
wire net1167;
wire net1168_c1;
wire net1168;
wire net1169_c1;
wire net1169;
wire net1170_c1;
wire net1170;
wire net1171_c1;
wire net1171;
wire net1172_c1;
wire net1172;
wire net1173_c1;
wire net1173;
wire net1174_c1;
wire net1174;
wire net1175_c1;
wire net1175;
wire net1176_c1;
wire net1176;
wire net1177_c1;
wire net1177;
wire net1178_c1;
wire net1178;
wire net1179_c1;
wire net1179;
wire net1180_c1;
wire net1180;
wire net1181_c1;
wire net1181;
wire net1182_c1;
wire net1182;
wire net1183_c1;
wire net1183;
wire net1184_c1;
wire net1184;
wire net1185_c1;
wire net1185;
wire net1186_c1;
wire net1186;
wire net1187_c1;
wire net1187;
wire net1188_c1;
wire net1188;
wire net1189_c1;
wire net1189;
wire net1190_c1;
wire net1190;
wire net1191_c1;
wire net1191;
wire net1192_c1;
wire net1192;
wire net1193_c1;
wire net1193;
wire net1194_c1;
wire net1194;
wire net1195_c1;
wire net1195;
wire net1196_c1;
wire net1196;
wire net1197_c1;
wire net1197;
wire net1198_c1;
wire net1198;
wire net1199_c1;
wire net1199;
wire net1200_c1;
wire net1200;
wire net1201_c1;
wire net1201;
wire net1202_c1;
wire net1202;
wire net1203_c1;
wire net1203;
wire net1204_c1;
wire net1204;
wire net1205_c1;
wire net1205;
wire net1206_c1;
wire net1206;
wire net1207_c1;
wire net1207;
wire net1208_c1;
wire net1208;
wire net1209_c1;
wire net1209;
wire net1210_c1;
wire net1210;
wire net1211_c1;
wire net1211;
wire GCLK_Pad;
wire net1212;
wire net1213_c1;
wire net1213;
wire net1214_c1;
wire net1214;
wire net1215_c1;
wire net1215;
wire net1216_c1;
wire net1216;
wire net1217_c1;
wire net1217;
wire net1218_c1;
wire net1218;
wire net1219_c1;
wire net1219;
wire net1220_c1;
wire net1220;
wire net1221_c1;
wire net1221;

DFFT DFFT_199__FPB_n658(net695,net58,net405_c1);
DFFT DFFT_105_state0_buf(net694,net194,net440_c1);
DFFT DFFT_251_state_obs1(net693,net370,net437_c1);
DFFT DFFT_245_state_obs0(net692,net324,net436_c1);
AND2T AND2T_100_n136(net691,net90,net430,net95_c1);
AND2T AND2T_110_n152(net690,net210,net195,net94_c1);
AND2T AND2T_107_n149(net689,net196,net169,net99_c1);
AND2T AND2T_108_n150(net688,net108,net432,net85_c1);
AND2T AND2T_109_n151(net687,net8,net434,net89_c1);
DFFT DFFT_101_state_obs0_buf(net686,net285,net281_c1);
DFFT DFFT_102_state_obs1_buf(net685,net286,net282_c1);
DFFT DFFT_103_state_obs2_buf(net684,net189,net283_c1);
DFFT DFFT_104_state_obs3_buf(net683,net280,net284_c1);
AND2T AND2T_8_n44(net682,net217,net279,net5_c1);
DFFT DFFT_106_state1_buf(net681,net201,net441_c1);
NOTT NOTT_9_n45(net680,net127,net8_c1);
XOR2T XOR2T_75_n111(net679,net206,net296,net61_c1);
AND2T AND2T_20_n56(net678,net112,net223,net20_c1);
AND2T AND2T_13_n49(net677,net193,net165,net26_c1);
AND2T AND2T_30_n66(net676,net247,net263,net30_c1);
AND2T AND2T_15_n51(net675,net104,net328,net2_c1);
AND2T AND2T_31_n67(net674,net132,net334,net35_c1);
AND2T AND2T_32_n68(net673,net215,net170,net40_c1);
AND2T AND2T_17_n53(net672,net11,net335,net7_c1);
AND2T AND2T_41_n77(net671,net150,net181,net43_c1);
AND2T AND2T_18_n54(net670,net1,net309,net11_c1);
AND2T AND2T_42_n78(net669,net251,net359,net47_c1);
AND2T AND2T_35_n71(net668,net227,net321,net13_c1);
AND2T AND2T_27_n63(net667,net220,net204,net14_c1);
AND2T AND2T_19_n55(net666,net259,net313,net15_c1);
AND2T AND2T_51_n87(net665,net230,net341,net49_c1);
AND2T AND2T_43_n79(net664,net145,net367,net50_c1);
AND2T AND2T_44_n80(net663,net233,net262,net17_c1);
AND2T AND2T_36_n72(net662,net116,net326,net18_c1);
AND2T AND2T_28_n64(net661,net232,net160,net19_c1);
AND2T AND2T_52_n88(net660,net126,net350,net52_c1);
AND2T AND2T_37_n73(net659,net237,net333,net23_c1);
AND2T AND2T_29_n65(net658,net133,net101,net24_c1);
AND2T AND2T_53_n89(net657,net149,net26,net54_c1);
AND2T AND2T_38_n74(net1082,net272,net342,net29_c1);
AND2T AND2T_62_n98(net656,net53,net358,net55_c1);
AND2T AND2T_55_n91(net655,net27,net374,net32_c1);
AND2T AND2T_39_n75(net654,net29,net254,net34_c1);
AND2T AND2T_63_n99(net653,net221,net183,net56_c1);
AND2T AND2T_48_n84(net652,net236,net274,net38_c1);
AND2T AND2T_49_n85(net651,net173,net1221,net42_c1);
AND2T AND2T_59_n95(net650,net45,net373,net48_c1);
DFFT DFFT_259_state_obs2(net649,net369,net438_c1);
DFFT DFFT_267_state_obs3(net648,net368,net439_c1);
DFFT DFFT_120__PIPL_n171(net647,net441,net286_c1);
OR2T OR2T_11_n47(net646,net12,net322,net16_c1);
OR2T OR2T_21_n57(net645,net250,net317,net25_c1);
OR2T OR2T_22_n58(net644,net7,net327,net31_c1);
OR2T OR2T_40_n76(net643,net34,net23,net39_c1);
OR2T OR2T_33_n69(net642,net40,net343,net44_c1);
OR2T OR2T_34_n70(net641,net44,net351,net9_c1);
OR2T OR2T_50_n86(net640,net42,net38,net46_c1);
OR2T OR2T_60_n96(net639,net143,net168,net51_c1);
OR2T OR2T_45_n81(net638,net224,net260,net22_c1);
OR2T OR2T_61_n97(net637,net140,net379,net53_c1);
OR2T OR2T_54_n90(net636,net54,net234,net27_c1);
OR2T OR2T_46_n82(net635,net22,net47,net28_c1);
OR2T OR2T_47_n83(net634,net28,net375,net33_c1);
OR2T OR2T_56_n92(net633,net32,net49,net37_c1);
OR2T OR2T_57_n93(net632,net37,net33,net41_c1);
OR2T OR2T_58_n94(net631,net41,net380,net45_c1);
DFFT DFFT_115__PIPL_n166(net630,net281,net287_c1);
DFFT DFFT_116__PIPL_n167(net629,net282,net288_c1);
NOTT NOTT_10_n46(net628,net255,net12_c1);
NOTT NOTT_12_n48(net627,net202,net21_c1);
NOTT NOTT_14_n50(net626,net257,net1_c1);
NOTT NOTT_23_n59(net625,net105,net36_c1);
NOTT NOTT_24_n60(net624,net267,net3_c1);
NOTT NOTT_16_n52(net623,net269,net4_c1);
NOTT NOTT_25_n61(net622,net192,net6_c1);
NOTT NOTT_26_n62(net621,net222,net10_c1);
DFFT DFFT_117__PIPL_n168(net620,net283,net289_c1);
DFFT DFFT_118__PIPL_n169(net619,net284,net290_c1);
DFFT DFFT_119__PIPL_n170(net618,net440,net285_c1);
AND2T AND2T_72_n108(net617,net76,net398,net80_c1);
AND2T AND2T_65_n101(net616,net243,net378,net58_c1);
AND2T AND2T_81_n117(net615,net276,net397,net83_c1);
AND2T AND2T_73_n109(net614,net158,net404,net84_c1);
AND2T AND2T_74_n110(net613,net213,net411,net59_c1);
AND2T AND2T_66_n102(net612,net130,net238,net60_c1);
AND2T AND2T_90_n126(net611,net82,net391,net87_c1);
AND2T AND2T_82_n118(net610,net83,net203,net88_c1);
AND2T AND2T_67_n103(net609,net248,net1219,net62_c1);
AND2T AND2T_91_n127(net608,net155,net410,net91_c1);
AND2T AND2T_76_n112(net824,net261,net416,net64_c1);
AND2T AND2T_92_n128(net607,net177,net1220,net96_c1);
AND2T AND2T_85_n121(net606,net208,net186,net66_c1);
AND2T AND2T_77_n113(net825,net199,net421,net67_c1);
AND2T AND2T_93_n129(net605,net114,net429,net98_c1);
AND2T AND2T_94_n130(net604,net73,net431,net69_c1);
AND2T AND2T_86_n122(net603,net66,net172,net70_c1);
AND2T AND2T_78_n114(net602,net268,net377,net71_c1);
DFFT DFFT_200__FPB_n659(net601,net137,net408_c1);
DFFT DFFT_121__FBL_n580(net600,net415,net291_c1);
DFFT DFFT_113__FPB_n164(net599,net129,net302_c1);
DFFT DFFT_201__FPB_n660(net598,net1218,net363_c1);
DFFT DFFT_122__FBL_n581(net597,net428,net292_c1);
DFFT DFFT_130__FBL_n589(net596,net312,net301_c1);
DFFT DFFT_114__FPB_n165(net595,net212,net303_c1);
DFFT DFFT_202__FPB_n661(net594,net363,net371_c1);
DFFT DFFT_210__FPB_n669(net593,net241,net421_c1);
DFFT DFFT_131__FBL_n590(net592,net316,net293_c1);
DFFT DFFT_123__FBL_n582(net591,net48,net294_c1);
DFFT DFFT_211__FPB_n670(net590,net148,net377_c1);
DFFT DFFT_203__FPB_n662(net589,net371,net376_c1);
DFFT DFFT_124__FBL_n583(net588,net256,net295_c1);
DFFT DFFT_212__FPB_n671(net587,net64,net386_c1);
DFFT DFFT_204__FPB_n663(net586,net376,net382_c1);
DFFT DFFT_132__FPB_n591(net585,net16,net385_c1);
DFFT DFFT_220__FPB_n679(net584,net424,net427_c1);
DFFT DFFT_140__FPB_n599(net583,net425,net428_c1);
DFFT DFFT_125__FBL_n584(net582,net304,net296_c1);
DFFT DFFT_141__FPB_n600(net581,net240,net304_c1);
DFFT DFFT_221__FPB_n680(net580,net427,net391_c1);
DFFT DFFT_213__FPB_n672(net579,net84,net392_c1);
DFFT DFFT_205__FPB_n664(net578,net382,net388_c1);
DFFT DFFT_133__FPB_n592(net577,net385,net390_c1);
DFFT DFFT_126__FBL_n585(net576,net305,net297_c1);
DFFT DFFT_142__FPB_n601(net575,net249,net305_c1);
DFFT DFFT_150__FPB_n609(net574,net190,net340_c1);
DFFT DFFT_222__FPB_n681(net573,net277,net394_c1);
DFFT DFFT_214__FPB_n673(net572,net205,net397_c1);
DFFT DFFT_206__FPB_n665(net571,net388,net398_c1);
DFFT DFFT_134__FPB_n593(net570,net390,net396_c1);
DFFT DFFT_230__FPB_n689(net569,net96,net433_c1);
DFFT DFFT_127__FBL_n586(net568,net167,net298_c1);
DFFT DFFT_151__FPB_n610(net567,net340,net306_c1);
DFFT DFFT_143__FPB_n602(net566,net146,net307_c1);
DFFT DFFT_231__FPB_n690(net565,net91,net402_c1);
DFFT DFFT_223__FPB_n682(net564,net1217,net400_c1);
DFFT DFFT_215__FPB_n674(net563,net70,net403_c1);
DFFT DFFT_207__FPB_n666(net562,net111,net404_c1);
DFFT DFFT_135__FPB_n594(net561,net396,net401_c1);
DFFT DFFT_128__FBL_n587(net560,net307,net299_c1);
OR2T OR2T_70_n106(net559,net68,net405,net72_c1);
OR2T OR2T_71_n107(net558,net72,net55,net76_c1);
OR2T OR2T_64_n100(net557,net56,net131,net57_c1);
OR2T OR2T_80_n116(net556,net1215,net392,net79_c1);
OR2T OR2T_83_n119(net555,net88,net163,net92_c1);
OR2T OR2T_84_n120(net554,net92,net139,net63_c1);
OR2T OR2T_68_n104(net553,net242,net393,net65_c1);
OR2T OR2T_69_n105(net552,net65,net399,net68_c1);
DFFT DFFT_152__FPB_n611(net551,net1216,net309_c1);
DFFT DFFT_144__FPB_n603(net550,net244,net308_c1);
DFFT DFFT_160__FPB_n619(net549,net184,net357_c1);
DFFT DFFT_232__FPB_n691(net548,net142,net406_c1);
DFFT DFFT_224__FPB_n683(net547,net400,net410_c1);
DFFT DFFT_216__FPB_n675(net546,net231,net407_c1);
DFFT DFFT_208__FPB_n667(net545,net110,net411_c1);
DFFT DFFT_136__FPB_n595(net544,net401,net409_c1);
OR2T OR2T_95_n131(net543,net214,net121,net73_c1);
OR2T OR2T_87_n123(net542,net239,net403,net74_c1);
OR2T OR2T_79_n115(net541,net71,net386,net75_c1);
DFFT DFFT_240__FPB_n699(net540,net287,net435_c1);
OR2T OR2T_96_n132(net539,net69,net98,net77_c1);
OR2T OR2T_88_n124(net538,net74,net63,net78_c1);
OR2T OR2T_97_n133(net537,net77,net252,net81_c1);
OR2T OR2T_89_n125(net536,net78,net79,net82_c1);
OR2T OR2T_98_n134(net535,net81,net433,net86_c1);
OR2T OR2T_99_n135(net534,net86,net402,net90_c1);
DFFT DFFT_129__FBL_n588(net533,net308,net300_c1);
DFFT DFFT_241__FPB_n700(net532,net435,net310_c1);
DFFT DFFT_161__FPB_n620(net531,net357,net311_c1);
DFFT DFFT_153__FPB_n612(net530,net115,net313_c1);
DFFT DFFT_145__FPB_n604(net529,net157,net312_c1);
DFFT DFFT_233__FPB_n692(net528,net406,net412_c1);
DFFT DFFT_225__FPB_n684(net527,net188,net413_c1);
DFFT DFFT_217__FPB_n676(net526,net407,net414_c1);
DFFT DFFT_209__FPB_n668(net525,net61,net416_c1);
DFFT DFFT_137__FPB_n596(net524,net409,net415_c1);
DFFT DFFT_242__FPB_n701(net523,net310,net314_c1);
DFFT DFFT_162__FPB_n621(net522,net311,net315_c1);
DFFT DFFT_154__FPB_n613(net521,net174,net317_c1);
DFFT DFFT_146__FPB_n605(net520,net153,net316_c1);
DFFT DFFT_250__FPB_n709(net519,net362,net370_c1);
DFFT DFFT_170__FPB_n629(net518,net154,net375_c1);
DFFT DFFT_234__FPB_n693(net517,net412,net417_c1);
DFFT DFFT_226__FPB_n685(net516,net413,net420_c1);
DFFT DFFT_218__FPB_n677(net515,net414,net418_c1);
DFFT DFFT_138__FPB_n597(net514,net31,net419_c1);
DFFT DFFT_243__FPB_n702(net513,net314,net318_c1);
DFFT DFFT_171__FPB_n630(net512,net159,net320_c1);
DFFT DFFT_163__FPB_n622(net511,net315,net321_c1);
DFFT DFFT_155__FPB_n614(net510,net25,net319_c1);
DFFT DFFT_147__FPB_n606(net509,net5,net322_c1);
DFFT DFFT_235__FPB_n694(net508,net417,net422_c1);
DFFT DFFT_227__FPB_n686(net507,net113,net423_c1);
DFFT DFFT_219__FPB_n678(net506,net418,net424_c1);
DFFT DFFT_139__FPB_n598(net505,net419,net425_c1);
DFFT DFFT_252__FPB_n711(net504,net289,net323_c1);
DFFT DFFT_244__FPB_n703(net503,net318,net324_c1);
DFFT DFFT_172__FPB_n631(net502,net271,net325_c1);
DFFT DFFT_164__FPB_n623(net501,net229,net326_c1);
DFFT DFFT_156__FPB_n615(net500,net319,net327_c1);
DFFT DFFT_148__FPB_n607(net499,net134,net328_c1);
DFFT DFFT_260__FPB_n719(net498,net290,net381_c1);
DFFT DFFT_180__FPB_n639(net497,net225,net384_c1);
DFFT DFFT_236__FPB_n695(net496,net422,net426_c1);
DFFT DFFT_228__FPB_n687(net495,net423,net429_c1);
DFFT DFFT_261__FPB_n720(net494,net381,net329_c1);
DFFT DFFT_253__FPB_n712(net493,net323,net330_c1);
DFFT DFFT_181__FPB_n640(net492,net384,net331_c1);
DFFT DFFT_173__FPB_n632(net491,net325,net332_c1);
DFFT DFFT_165__FPB_n624(net490,net266,net333_c1);
DFFT DFFT_157__FPB_n616(net489,net103,net334_c1);
DFFT DFFT_149__FPB_n608(net488,net4,net335_c1);
DFFT DFFT_237__FPB_n696(net487,net1214,net430_c1);
DFFT DFFT_229__FPB_n688(net486,net207,net431_c1);
DFFT DFFT_262__FPB_n721(net1210,net329,net336_c1);
DFFT DFFT_254__FPB_n713(net485,net330,net337_c1);
DFFT DFFT_246__FPB_n705(net484,net288,net338_c1);
DFFT DFFT_182__FPB_n641(net483,net331,net339_c1);
DFFT DFFT_174__FPB_n633(net482,net332,net341_c1);
DFFT DFFT_166__FPB_n625(net1083,net138,net342_c1);
DFFT DFFT_158__FPB_n617(net481,net30,net343_c1);
DFFT DFFT_190__FPB_n649(net480,net389,net395_c1);
DFFT DFFT_238__FPB_n697(net479,net102,net432_c1);
SPLITT Split_300_n759(net50,net168_c1,net260_c1);
SPLITT Split_301_n760(net17,net131_c1,net224_c1);
SPLITT Split_302_n761(net46,net139_c1,net230_c1);
SPLITT Split_310_n769(net67,net177_c1,net268_c1);
SPLITT Split_303_n762(net52,net143_c1,net234_c1);
SPLITT Split_311_n770(net87,net141_c1,net235_c1);
SPLITT Split_304_n763(net51,net147_c1,net239_c1);
SPLITT Split_312_n771(net235,net146_c1,net240_c1);
SPLITT Split_320_n779(net175,net183_c1,net274_c1);
SPLITT Split_305_n764(net57,net155_c1,net243_c1);
SPLITT Split_313_n772(net141,net153_c1,net244_c1);
SPLITT Split_321_n780(net89,net151_c1,net245_c1);
SPLITT Split_306_n765(net60,net158_c1,net248_c1);
SPLITT Split_314_n773(net95,net157_c1,net249_c1);
SPLITT Split_322_n781(net245,net160_c1,net250_c1);
SPLITT Split_330_n789(net93,net187_c1,net278_c1);
SPLITT Split_307_n766(net62,net162_c1,net252_c1);
SPLITT Split_315_n774(net99,net161_c1,net253_c1);
SPLITT Split_323_n782(net151,net164_c1,net254_c1);
SPLITT Split_331_n790(net278,net165_c1,net255_c1);
SPLITT Split_308_n767(net80,net167_c1,net256_c1);
SPLITT Split_316_n775(net253,net170_c1,net257_c1);
SPLITT Split_324_n783(net94,net166_c1,net258_c1);
SPLITT Split_332_n791(net187,net169_c1,net259_c1);
SPLITT Split_340_n799(net292,net190_c1,net280_c1);
SPLITT Split_341_n800(net294,net100_c1,net191_c1);
SPLITT Split_309_n768(net59,net172_c1,net261_c1);
SPLITT Split_317_n776(net161,net173_c1,net262_c1);
SPLITT Split_325_n784(net258,net174_c1,net263_c1);
SPLITT Split_333_n792(net302,net171_c1,net264_c1);
SPLITT Split_342_n801(net191,net101_c1,net192_c1);
SPLITT Split_270_n729(net21,net136_c1,net228_c1);
SPLITT Split_350_n809(net122,net138_c1,net229_c1);
SPLITT Split_318_n777(net85,net175_c1,net265_c1);
SPLITT Split_326_n785(net166,net176_c1,net266_c1);
SPLITT Split_334_n793(net264,net178_c1,net267_c1);
SPLITT Split_271_n730(net228,net104_c1,net193_c1);
SPLITT Split_343_n802(net100,net103_c1,net194_c1);
SPLITT Split_351_n810(net299,net102_c1,net195_c1);
SPLITT Split_319_n778(net265,net181_c1,net269_c1);
SPLITT Split_327_n786(net97,net179_c1,net270_c1);
SPLITT Split_335_n794(net171,net180_c1,net271_c1);
SPLITT Split_272_n731(net136,net108_c1,net196_c1);
SPLITT Split_344_n803(net295,net107_c1,net197_c1);
SPLITT Split_352_n811(net301,net106_c1,net198_c1);
SPLITT Split_280_n739(net3,net148_c1,net238_c1);
SPLITT Split_328_n787(net270,net184_c1,net272_c1);
SPLITT Split_336_n795(net303,net182_c1,net273_c1);
SPLITT Split_273_n732(net2,net111_c1,net199_c1);
SPLITT Split_281_n740(net6,net109_c1,net200_c1);
SPLITT Split_345_n804(net197,net110_c1,net201_c1);
SPLITT Split_353_n812(net198,net112_c1,net202_c1);
SPLITT Split_329_n788(net179,net185_c1,net275_c1);
SPLITT Split_337_n796(net273,net186_c1,net276_c1);
DFFT DFFT_263__FPB_n722(net1211,net336,net344_c1);
DFFT DFFT_255__FPB_n714(net478,net337,net345_c1);
DFFT DFFT_247__FPB_n706(net477,net338,net346_c1);
DFFT DFFT_191__FPB_n650(net476,net395,net347_c1);
DFFT DFFT_183__FPB_n642(net475,net339,net348_c1);
DFFT DFFT_175__FPB_n634(net474,net125,net350_c1);
DFFT DFFT_167__FPB_n626(net473,net178,net349_c1);
DFFT DFFT_159__FPB_n618(net472,net19,net351_c1);
SPLITT Split_274_n733(net15,net114_c1,net203_c1);
SPLITT Split_282_n741(net200,net116_c1,net204_c1);
SPLITT Split_346_n805(net107,net113_c1,net205_c1);
SPLITT Split_354_n813(net106,net115_c1,net206_c1);
SPLITT Split_290_n749(net152,net159_c1,net247_c1);
DFFT DFFT_239__FPB_n698(net471,net120,net434_c1);
SPLITT Split_338_n797(net182,net188_c1,net277_c1);
SPLITT Split_275_n734(net20,net119_c1,net207_c1);
SPLITT Split_283_n742(net109,net121_c1,net208_c1);
SPLITT Split_291_n750(net35,net118_c1,net209_c1);
SPLITT Split_347_n806(net297,net120_c1,net210_c1);
SPLITT Split_355_n814(net293,net117_c1,net211_c1);
SPLITT Split_339_n798(net291,net189_c1,net279_c1);
SPLITT Split_268_n727(net0,net123_c1,net212_c1);
SPLITT Split_276_n735(net119,net125_c1,net213_c1);
SPLITT Split_284_n743(net10,net124_c1,net214_c1);
SPLITT Split_292_n751(net209,net126_c1,net215_c1);
SPLITT Split_348_n807(net298,net122_c1,net216_c1);
SPLITT Split_356_n815(net211,net127_c1,net217_c1);
SPLITT Split_269_n728(net123,net129_c1,net218_c1);
SPLITT Split_277_n736(net36,net128_c1,net219_c1);
SPLITT Split_285_n744(net124,net132_c1,net220_c1);
SPLITT Split_293_n752(net118,net130_c1,net221_c1);
SPLITT Split_349_n808(net216,net133_c1,net222_c1);
SPLITT Split_357_n816(net117,net134_c1,net223_c1);
SPLITT Split_278_n737(net219,net137_c1,net225_c1);
SPLITT Split_286_n745(net14,net135_c1,net226_c1);
SPLITT Split_294_n753(net9,net140_c1,net227_c1);
SPLITT Split_279_n738(net128,net142_c1,net231_c1);
SPLITT Split_287_n746(net226,net145_c1,net232_c1);
SPLITT Split_295_n754(net18,net144_c1,net233_c1);
SPLITT Split_288_n747(net135,net149_c1,net236_c1);
SPLITT Split_296_n755(net144,net150_c1,net237_c1);
SPLITT Split_289_n748(net24,net152_c1,net241_c1);
SPLITT Split_297_n756(net39,net154_c1,net242_c1);
SPLITT Split_298_n757(net43,net156_c1,net246_c1);
SPLITT Split_299_n758(net156,net163_c1,net251_c1);
NOTT NOTT_111_n153(net470,net218,net97_c1);
NOTT NOTT_112_n160(net469,net300,net93_c1);
DFFT DFFT_264__FPB_n723(net468,net344,net352_c1);
DFFT DFFT_256__FPB_n715(net952,net345,net353_c1);
DFFT DFFT_248__FPB_n707(net467,net346,net354_c1);
DFFT DFFT_192__FPB_n651(net466,net347,net358_c1);
DFFT DFFT_184__FPB_n643(net465,net348,net355_c1);
DFFT DFFT_176__FPB_n635(net464,net275,net356_c1);
DFFT DFFT_168__FPB_n627(net463,net349,net359_c1);
DFFT DFFT_265__FPB_n724(net462,net352,net360_c1);
DFFT DFFT_257__FPB_n716(net953,net353,net361_c1);
DFFT DFFT_249__FPB_n708(net461,net354,net362_c1);
DFFT DFFT_193__FPB_n652(net460,net185,net364_c1);
DFFT DFFT_185__FPB_n644(net459,net355,net365_c1);
DFFT DFFT_177__FPB_n636(net458,net356,net366_c1);
DFFT DFFT_169__FPB_n628(net457,net176,net367_c1);
DFFT DFFT_266__FPB_n725(net456,net360,net368_c1);
DFFT DFFT_258__FPB_n717(net455,net361,net369_c1);
DFFT DFFT_194__FPB_n653(net454,net364,net372_c1);
DFFT DFFT_186__FPB_n645(net453,net365,net373_c1);
DFFT DFFT_178__FPB_n637(net452,net366,net374_c1);
DFFT DFFT_195__FPB_n654(net451,net372,net378_c1);
DFFT DFFT_187__FPB_n646(net450,net147,net379_c1);
DFFT DFFT_179__FPB_n638(net449,net13,net380_c1);
DFFT DFFT_196__FPB_n655(net448,net164,net387_c1);
DFFT DFFT_188__FPB_n647(net447,net180,net383_c1);
DFFT DFFT_197__FPB_n656(net446,net246,net393_c1);
DFFT DFFT_189__FPB_n648(net445,net1213,net389_c1);
DFFT DFFT_198__FPB_n657(net444,net162,net399_c1);
SPLITT SplitCLK_0_261(net1209,net1210_c1,net1211_c1);
SPLITT SplitCLK_0_262(net1204,net1209_c1,net1208_c1);
SPLITT SplitCLK_6_263(net1205,net1207_c1,net1206_c1);
SPLITT SplitCLK_0_264(net1196,net1205_c1,net1204_c1);
SPLITT SplitCLK_0_265(net1198,net1203_c1,net1202_c1);
SPLITT SplitCLK_2_266(net1199,net1200_c1,net1201_c1);
SPLITT SplitCLK_6_267(net1197,net1198_c1,net1199_c1);
SPLITT SplitCLK_4_268(net1180,net1197_c1,net1196_c1);
SPLITT SplitCLK_0_269(net1190,net1194_c1,net1195_c1);
SPLITT SplitCLK_6_270(net1191,net1192_c1,net1193_c1);
SPLITT SplitCLK_6_271(net1182,net1190_c1,net1191_c1);
SPLITT SplitCLK_0_272(net1184,net1188_c1,net1189_c1);
SPLITT SplitCLK_2_273(net1185,net1186_c1,net1187_c1);
SPLITT SplitCLK_4_274(net1183,net1185_c1,net1184_c1);
SPLITT SplitCLK_2_275(net1181,net1183_c1,net1182_c1);
SPLITT SplitCLK_6_276(net1148,net1180_c1,net1181_c1);
SPLITT SplitCLK_0_277(net1174,net1179_c1,net1178_c1);
SPLITT SplitCLK_2_278(net1175,net1176_c1,net1177_c1);
SPLITT SplitCLK_4_279(net1166,net1175_c1,net1174_c1);
SPLITT SplitCLK_0_280(net1168,net1172_c1,net1173_c1);
SPLITT SplitCLK_0_281(net1169,net1170_c1,net1171_c1);
SPLITT SplitCLK_4_282(net1167,net1169_c1,net1168_c1);
SPLITT SplitCLK_0_283(net1150,net1166_c1,net1167_c1);
SPLITT SplitCLK_0_284(net1160,net1164_c1,net1165_c1);
SPLITT SplitCLK_4_285(net1161,net1162_c1,net1163_c1);
SPLITT SplitCLK_6_286(net1152,net1160_c1,net1161_c1);
SPLITT SplitCLK_0_287(net1154,net1159_c1,net1158_c1);
SPLITT SplitCLK_2_288(net1155,net1156_c1,net1157_c1);
SPLITT SplitCLK_4_289(net1153,net1155_c1,net1154_c1);
SPLITT SplitCLK_2_290(net1151,net1153_c1,net1152_c1);
SPLITT SplitCLK_4_291(net1149,net1151_c1,net1150_c1);
SPLITT SplitCLK_0_292(net1084,net1148_c1,net1149_c1);
SPLITT SplitCLK_4_293(net1142,net1146_c1,net1147_c1);
SPLITT SplitCLK_6_294(net1143,net1144_c1,net1145_c1);
SPLITT SplitCLK_6_295(net1134,net1142_c1,net1143_c1);
SPLITT SplitCLK_4_296(net1136,net1140_c1,net1141_c1);
SPLITT SplitCLK_4_297(net1137,net1139_c1,net1138_c1);
SPLITT SplitCLK_0_298(net1135,net1136_c1,net1137_c1);
SPLITT SplitCLK_4_299(net1118,net1135_c1,net1134_c1);
SPLITT SplitCLK_0_300(net1128,net1133_c1,net1132_c1);
SPLITT SplitCLK_6_301(net1129,net1131_c1,net1130_c1);
SPLITT SplitCLK_2_302(net1120,net1128_c1,net1129_c1);
SPLITT SplitCLK_0_303(net1122,net1126_c1,net1127_c1);
SPLITT SplitCLK_2_304(net1123,net1124_c1,net1125_c1);
SPLITT SplitCLK_4_305(net1121,net1123_c1,net1122_c1);
SPLITT SplitCLK_6_306(net1119,net1121_c1,net1120_c1);
SPLITT SplitCLK_2_307(net1086,net1118_c1,net1119_c1);
SPLITT SplitCLK_0_308(net1112,net1116_c1,net1117_c1);
SPLITT SplitCLK_6_309(net1113,net1114_c1,net1115_c1);
SPLITT SplitCLK_6_310(net1104,net1112_c1,net1113_c1);
SPLITT SplitCLK_4_311(net1106,net1110_c1,net1111_c1);
SPLITT SplitCLK_6_312(net1107,net1108_c1,net1109_c1);
SPLITT SplitCLK_4_313(net1105,net1107_c1,net1106_c1);
SPLITT SplitCLK_0_314(net1088,net1104_c1,net1105_c1);
SPLITT SplitCLK_4_315(net1098,net1103_c1,net1102_c1);
SPLITT SplitCLK_6_316(net1099,net1100_c1,net1101_c1);
SPLITT SplitCLK_6_317(net1090,net1098_c1,net1099_c1);
SPLITT SplitCLK_4_318(net1092,net1096_c1,net1097_c1);
SPLITT SplitCLK_2_319(net1093,net1094_c1,net1095_c1);
SPLITT SplitCLK_4_320(net1091,net1093_c1,net1092_c1);
SPLITT SplitCLK_2_321(net1089,net1091_c1,net1090_c1);
SPLITT SplitCLK_4_322(net1087,net1089_c1,net1088_c1);
SPLITT SplitCLK_2_323(net1085,net1087_c1,net1086_c1);
SPLITT SplitCLK_6_324(net954,net1084_c1,net1085_c1);
SPLITT SplitCLK_4_325(net1081,net1083_c1,net1082_c1);
SPLITT SplitCLK_2_326(net1076,net1080_c1,net1081_c1);
SPLITT SplitCLK_6_327(net1077,net1079_c1,net1078_c1);
SPLITT SplitCLK_0_328(net1068,net1077_c1,net1076_c1);
SPLITT SplitCLK_0_329(net1070,net1075_c1,net1074_c1);
SPLITT SplitCLK_2_330(net1071,net1073_c1,net1072_c1);
SPLITT SplitCLK_4_331(net1069,net1071_c1,net1070_c1);
SPLITT SplitCLK_4_332(net1052,net1068_c1,net1069_c1);
SPLITT SplitCLK_0_333(net1062,net1066_c1,net1067_c1);
SPLITT SplitCLK_6_334(net1063,net1065_c1,net1064_c1);
SPLITT SplitCLK_6_335(net1054,net1062_c1,net1063_c1);
SPLITT SplitCLK_4_336(net1056,net1060_c1,net1061_c1);
SPLITT SplitCLK_2_337(net1057,net1058_c1,net1059_c1);
SPLITT SplitCLK_4_338(net1055,net1057_c1,net1056_c1);
SPLITT SplitCLK_6_339(net1053,net1055_c1,net1054_c1);
SPLITT SplitCLK_6_340(net1020,net1052_c1,net1053_c1);
SPLITT SplitCLK_4_341(net1046,net1050_c1,net1051_c1);
SPLITT SplitCLK_6_342(net1047,net1049_c1,net1048_c1);
SPLITT SplitCLK_4_343(net1038,net1047_c1,net1046_c1);
SPLITT SplitCLK_0_344(net1040,net1045_c1,net1044_c1);
SPLITT SplitCLK_4_345(net1041,net1042_c1,net1043_c1);
SPLITT SplitCLK_4_346(net1039,net1041_c1,net1040_c1);
SPLITT SplitCLK_0_347(net1022,net1038_c1,net1039_c1);
SPLITT SplitCLK_0_348(net1032,net1037_c1,net1036_c1);
SPLITT SplitCLK_6_349(net1033,net1034_c1,net1035_c1);
SPLITT SplitCLK_6_350(net1024,net1032_c1,net1033_c1);
SPLITT SplitCLK_4_351(net1026,net1030_c1,net1031_c1);
SPLITT SplitCLK_2_352(net1027,net1028_c1,net1029_c1);
SPLITT SplitCLK_4_353(net1025,net1027_c1,net1026_c1);
SPLITT SplitCLK_4_354(net1023,net1024_c1,net1025_c1);
SPLITT SplitCLK_4_355(net1021,net1023_c1,net1022_c1);
SPLITT SplitCLK_4_356(net956,net1021_c1,net1020_c1);
SPLITT SplitCLK_0_357(net1014,net1018_c1,net1019_c1);
SPLITT SplitCLK_6_358(net1015,net1016_c1,net1017_c1);
SPLITT SplitCLK_4_359(net1006,net1015_c1,net1014_c1);
SPLITT SplitCLK_0_360(net1008,net1013_c1,net1012_c1);
SPLITT SplitCLK_2_361(net1009,net1011_c1,net1010_c1);
SPLITT SplitCLK_4_362(net1007,net1009_c1,net1008_c1);
SPLITT SplitCLK_0_363(net990,net1006_c1,net1007_c1);
SPLITT SplitCLK_0_364(net1000,net1005_c1,net1004_c1);
SPLITT SplitCLK_6_365(net1001,net1002_c1,net1003_c1);
SPLITT SplitCLK_4_366(net992,net1001_c1,net1000_c1);
SPLITT SplitCLK_4_367(net994,net999_c1,net998_c1);
SPLITT SplitCLK_0_368(net995,net996_c1,net997_c1);
SPLITT SplitCLK_4_369(net993,net995_c1,net994_c1);
SPLITT SplitCLK_2_370(net991,net993_c1,net992_c1);
SPLITT SplitCLK_6_371(net958,net990_c1,net991_c1);
SPLITT SplitCLK_0_372(net984,net988_c1,net989_c1);
SPLITT SplitCLK_6_373(net985,net987_c1,net986_c1);
SPLITT SplitCLK_2_374(net976,net984_c1,net985_c1);
SPLITT SplitCLK_0_375(net978,net982_c1,net983_c1);
SPLITT SplitCLK_4_376(net979,net980_c1,net981_c1);
SPLITT SplitCLK_4_377(net977,net979_c1,net978_c1);
SPLITT SplitCLK_0_378(net960,net976_c1,net977_c1);
SPLITT SplitCLK_0_379(net970,net975_c1,net974_c1);
SPLITT SplitCLK_4_380(net971,net973_c1,net972_c1);
SPLITT SplitCLK_2_381(net962,net970_c1,net971_c1);
SPLITT SplitCLK_0_382(net964,net969_c1,net968_c1);
SPLITT SplitCLK_2_383(net965,net966_c1,net967_c1);
SPLITT SplitCLK_2_384(net963,net964_c1,net965_c1);
SPLITT SplitCLK_4_385(net961,net963_c1,net962_c1);
SPLITT SplitCLK_4_386(net959,net961_c1,net960_c1);
SPLITT SplitCLK_2_387(net957,net959_c1,net958_c1);
SPLITT SplitCLK_4_388(net955,net957_c1,net956_c1);
SPLITT SplitCLK_0_389(net442,net954_c1,net955_c1);
SPLITT SplitCLK_0_390(net951,net952_c1,net953_c1);
SPLITT SplitCLK_0_391(net946,net951_c1,net950_c1);
SPLITT SplitCLK_2_392(net947,net948_c1,net949_c1);
SPLITT SplitCLK_0_393(net938,net947_c1,net946_c1);
SPLITT SplitCLK_4_394(net940,net944_c1,net945_c1);
SPLITT SplitCLK_6_395(net941,net942_c1,net943_c1);
SPLITT SplitCLK_4_396(net939,net941_c1,net940_c1);
SPLITT SplitCLK_4_397(net922,net938_c1,net939_c1);
SPLITT SplitCLK_0_398(net932,net937_c1,net936_c1);
SPLITT SplitCLK_6_399(net933,net935_c1,net934_c1);
SPLITT SplitCLK_0_400(net924,net933_c1,net932_c1);
SPLITT SplitCLK_0_401(net926,net931_c1,net930_c1);
SPLITT SplitCLK_6_402(net927,net928_c1,net929_c1);
SPLITT SplitCLK_2_403(net925,net926_c1,net927_c1);
SPLITT SplitCLK_2_404(net923,net925_c1,net924_c1);
SPLITT SplitCLK_6_405(net890,net922_c1,net923_c1);
SPLITT SplitCLK_0_406(net916,net921_c1,net920_c1);
SPLITT SplitCLK_2_407(net917,net918_c1,net919_c1);
SPLITT SplitCLK_6_408(net908,net916_c1,net917_c1);
SPLITT SplitCLK_0_409(net910,net915_c1,net914_c1);
SPLITT SplitCLK_4_410(net911,net913_c1,net912_c1);
SPLITT SplitCLK_4_411(net909,net911_c1,net910_c1);
SPLITT SplitCLK_0_412(net892,net908_c1,net909_c1);
SPLITT SplitCLK_0_413(net902,net906_c1,net907_c1);
SPLITT SplitCLK_2_414(net903,net905_c1,net904_c1);
SPLITT SplitCLK_0_415(net894,net903_c1,net902_c1);
SPLITT SplitCLK_0_416(net896,net901_c1,net900_c1);
SPLITT SplitCLK_6_417(net897,net899_c1,net898_c1);
SPLITT SplitCLK_2_418(net895,net896_c1,net897_c1);
SPLITT SplitCLK_4_419(net893,net895_c1,net894_c1);
SPLITT SplitCLK_4_420(net891,net893_c1,net892_c1);
SPLITT SplitCLK_0_421(net826,net890_c1,net891_c1);
SPLITT SplitCLK_0_422(net884,net889_c1,net888_c1);
SPLITT SplitCLK_6_423(net885,net887_c1,net886_c1);
SPLITT SplitCLK_0_424(net876,net885_c1,net884_c1);
SPLITT SplitCLK_0_425(net878,net882_c1,net883_c1);
SPLITT SplitCLK_6_426(net879,net880_c1,net881_c1);
SPLITT SplitCLK_4_427(net877,net879_c1,net878_c1);
SPLITT SplitCLK_4_428(net860,net876_c1,net877_c1);
SPLITT SplitCLK_0_429(net870,net875_c1,net874_c1);
SPLITT SplitCLK_6_430(net871,net873_c1,net872_c1);
SPLITT SplitCLK_6_431(net862,net870_c1,net871_c1);
SPLITT SplitCLK_4_432(net864,net869_c1,net868_c1);
SPLITT SplitCLK_6_433(net865,net866_c1,net867_c1);
SPLITT SplitCLK_4_434(net863,net865_c1,net864_c1);
SPLITT SplitCLK_2_435(net861,net863_c1,net862_c1);
SPLITT SplitCLK_6_436(net828,net860_c1,net861_c1);
SPLITT SplitCLK_0_437(net854,net858_c1,net859_c1);
SPLITT SplitCLK_2_438(net855,net856_c1,net857_c1);
SPLITT SplitCLK_2_439(net846,net854_c1,net855_c1);
SPLITT SplitCLK_4_440(net848,net853_c1,net852_c1);
SPLITT SplitCLK_6_441(net849,net850_c1,net851_c1);
SPLITT SplitCLK_2_442(net847,net848_c1,net849_c1);
SPLITT SplitCLK_4_443(net830,net847_c1,net846_c1);
SPLITT SplitCLK_4_444(net840,net845_c1,net844_c1);
SPLITT SplitCLK_2_445(net841,net842_c1,net843_c1);
SPLITT SplitCLK_6_446(net832,net840_c1,net841_c1);
SPLITT SplitCLK_4_447(net834,net839_c1,net838_c1);
SPLITT SplitCLK_0_448(net835,net836_c1,net837_c1);
SPLITT SplitCLK_4_449(net833,net835_c1,net834_c1);
SPLITT SplitCLK_2_450(net831,net833_c1,net832_c1);
SPLITT SplitCLK_4_451(net829,net831_c1,net830_c1);
SPLITT SplitCLK_2_452(net827,net829_c1,net828_c1);
SPLITT SplitCLK_6_453(net696,net826_c1,net827_c1);
SPLITT SplitCLK_0_454(net823,net824_c1,net825_c1);
SPLITT SplitCLK_0_455(net818,net823_c1,net822_c1);
SPLITT SplitCLK_6_456(net819,net821_c1,net820_c1);
SPLITT SplitCLK_2_457(net810,net818_c1,net819_c1);
SPLITT SplitCLK_0_458(net812,net816_c1,net817_c1);
SPLITT SplitCLK_2_459(net813,net815_c1,net814_c1);
SPLITT SplitCLK_4_460(net811,net813_c1,net812_c1);
SPLITT SplitCLK_4_461(net794,net810_c1,net811_c1);
SPLITT SplitCLK_0_462(net804,net809_c1,net808_c1);
SPLITT SplitCLK_4_463(net805,net806_c1,net807_c1);
SPLITT SplitCLK_2_464(net796,net804_c1,net805_c1);
SPLITT SplitCLK_4_465(net798,net803_c1,net802_c1);
SPLITT SplitCLK_2_466(net799,net801_c1,net800_c1);
SPLITT SplitCLK_4_467(net797,net799_c1,net798_c1);
SPLITT SplitCLK_2_468(net795,net797_c1,net796_c1);
SPLITT SplitCLK_6_469(net762,net794_c1,net795_c1);
SPLITT SplitCLK_4_470(net788,net793_c1,net792_c1);
SPLITT SplitCLK_6_471(net789,net791_c1,net790_c1);
SPLITT SplitCLK_6_472(net780,net788_c1,net789_c1);
SPLITT SplitCLK_0_473(net782,net787_c1,net786_c1);
SPLITT SplitCLK_6_474(net783,net785_c1,net784_c1);
SPLITT SplitCLK_4_475(net781,net783_c1,net782_c1);
SPLITT SplitCLK_4_476(net764,net780_c1,net781_c1);
SPLITT SplitCLK_0_477(net774,net778_c1,net779_c1);
SPLITT SplitCLK_2_478(net775,net776_c1,net777_c1);
SPLITT SplitCLK_6_479(net766,net774_c1,net775_c1);
SPLITT SplitCLK_0_480(net768,net772_c1,net773_c1);
SPLITT SplitCLK_6_481(net769,net771_c1,net770_c1);
SPLITT SplitCLK_4_482(net767,net769_c1,net768_c1);
SPLITT SplitCLK_2_483(net765,net767_c1,net766_c1);
SPLITT SplitCLK_4_484(net763,net765_c1,net764_c1);
SPLITT SplitCLK_0_485(net698,net762_c1,net763_c1);
SPLITT SplitCLK_0_486(net756,net760_c1,net761_c1);
SPLITT SplitCLK_6_487(net757,net759_c1,net758_c1);
SPLITT SplitCLK_6_488(net748,net756_c1,net757_c1);
SPLITT SplitCLK_0_489(net750,net755_c1,net754_c1);
SPLITT SplitCLK_2_490(net751,net752_c1,net753_c1);
SPLITT SplitCLK_4_491(net749,net751_c1,net750_c1);
SPLITT SplitCLK_0_492(net732,net748_c1,net749_c1);
SPLITT SplitCLK_0_493(net742,net746_c1,net747_c1);
SPLITT SplitCLK_4_494(net743,net745_c1,net744_c1);
SPLITT SplitCLK_2_495(net734,net743_c1,net742_c1);
SPLITT SplitCLK_0_496(net736,net740_c1,net741_c1);
SPLITT SplitCLK_6_497(net737,net738_c1,net739_c1);
SPLITT SplitCLK_4_498(net735,net737_c1,net736_c1);
SPLITT SplitCLK_2_499(net733,net735_c1,net734_c1);
SPLITT SplitCLK_6_500(net700,net732_c1,net733_c1);
SPLITT SplitCLK_0_501(net726,net731_c1,net730_c1);
SPLITT SplitCLK_6_502(net727,net728_c1,net729_c1);
SPLITT SplitCLK_4_503(net718,net727_c1,net726_c1);
SPLITT SplitCLK_4_504(net720,net725_c1,net724_c1);
SPLITT SplitCLK_2_505(net721,net723_c1,net722_c1);
SPLITT SplitCLK_4_506(net719,net721_c1,net720_c1);
SPLITT SplitCLK_4_507(net702,net719_c1,net718_c1);
SPLITT SplitCLK_0_508(net712,net717_c1,net716_c1);
SPLITT SplitCLK_2_509(net713,net715_c1,net714_c1);
SPLITT SplitCLK_6_510(net704,net712_c1,net713_c1);
SPLITT SplitCLK_4_511(net706,net711_c1,net710_c1);
SPLITT SplitCLK_6_512(net707,net708_c1,net709_c1);
SPLITT SplitCLK_4_513(net705,net707_c1,net706_c1);
SPLITT SplitCLK_2_514(net703,net705_c1,net704_c1);
SPLITT SplitCLK_4_515(net701,net703_c1,net702_c1);
SPLITT SplitCLK_4_516(net699,net700_c1,net701_c1);
SPLITT SplitCLK_4_517(net697,net699_c1,net698_c1);
SPLITT SplitCLK_2_518(net443,net697_c1,net696_c1);
wire dummy0;
SPLITT SplitCLK_2_519(net986,net695_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_4_520(net888,net694_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_521(net889,net693_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_522(net872,net692_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_4_523(net778,net691_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_2_524(net1162,net690_c1,dummy5);
wire dummy6;
SPLITT SplitCLK_2_525(net1102,net689_c1,dummy6);
wire dummy7;
SPLITT SplitCLK_2_526(net1103,net688_c1,dummy7);
wire dummy8;
SPLITT SplitCLK_4_527(net1202,net687_c1,dummy8);
wire dummy9;
SPLITT SplitCLK_2_528(net880,net686_c1,dummy9);
wire dummy10;
SPLITT SplitCLK_4_529(net936,net685_c1,dummy10);
wire dummy11;
SPLITT SplitCLK_2_530(net1126,net684_c1,dummy11);
wire dummy12;
SPLITT SplitCLK_2_531(net1194,net683_c1,dummy12);
wire dummy13;
SPLITT SplitCLK_4_532(net1124,net682_c1,dummy13);
wire dummy14;
SPLITT SplitCLK_4_533(net930,net681_c1,dummy14);
wire dummy15;
SPLITT SplitCLK_4_534(net1200,net680_c1,dummy15);
wire dummy16;
SPLITT SplitCLK_2_535(net906,net679_c1,dummy16);
wire dummy17;
SPLITT SplitCLK_2_536(net904,net678_c1,dummy17);
wire dummy18;
SPLITT SplitCLK_2_537(net1100,net677_c1,dummy18);
wire dummy19;
SPLITT SplitCLK_2_538(net912,net676_c1,dummy19);
wire dummy20;
SPLITT SplitCLK_4_539(net920,net675_c1,dummy20);
wire dummy21;
SPLITT SplitCLK_2_540(net913,net674_c1,dummy21);
wire dummy22;
SPLITT SplitCLK_4_541(net905,net673_c1,dummy22);
wire dummy23;
SPLITT SplitCLK_2_542(net1140,net672_c1,dummy23);
wire dummy24;
SPLITT SplitCLK_4_543(net1158,net671_c1,dummy24);
wire dummy25;
SPLITT SplitCLK_4_544(net1141,net670_c1,dummy25);
wire dummy26;
SPLITT SplitCLK_2_545(net814,net669_c1,dummy26);
wire dummy27;
SPLITT SplitCLK_4_546(net1074,net668_c1,dummy27);
wire dummy28;
SPLITT SplitCLK_4_547(net1094,net667_c1,dummy28);
wire dummy29;
SPLITT SplitCLK_2_548(net898,net666_c1,dummy29);
wire dummy30;
SPLITT SplitCLK_2_549(net988,net665_c1,dummy30);
wire dummy31;
SPLITT SplitCLK_2_550(net1172,net664_c1,dummy31);
wire dummy32;
SPLITT SplitCLK_2_551(net1156,net663_c1,dummy32);
wire dummy33;
SPLITT SplitCLK_4_552(net1173,net662_c1,dummy33);
wire dummy34;
SPLITT SplitCLK_2_553(net1101,net661_c1,dummy34);
wire dummy35;
SPLITT SplitCLK_4_554(net914,net660_c1,dummy35);
wire dummy36;
SPLITT SplitCLK_4_555(net1170,net659_c1,dummy36);
wire dummy37;
SPLITT SplitCLK_2_556(net758,net658_c1,dummy37);
wire dummy38;
SPLITT SplitCLK_4_557(net1159,net657_c1,dummy38);
wire dummy39;
SPLITT SplitCLK_4_558(net792,net656_c1,dummy39);
wire dummy40;
SPLITT SplitCLK_4_559(net1058,net655_c1,dummy40);
wire dummy41;
SPLITT SplitCLK_2_560(net1080,net654_c1,dummy41);
wire dummy42;
SPLITT SplitCLK_4_561(net1110,net653_c1,dummy42);
wire dummy43;
SPLITT SplitCLK_2_562(net1157,net652_c1,dummy43);
wire dummy44;
SPLITT SplitCLK_2_563(net1096,net651_c1,dummy44);
wire dummy45;
SPLITT SplitCLK_4_564(net738,net650_c1,dummy45);
wire dummy46;
SPLITT SplitCLK_2_565(net937,net649_c1,dummy46);
wire dummy47;
SPLITT SplitCLK_2_566(net1130,net648_c1,dummy47);
wire dummy48;
SPLITT SplitCLK_2_567(net931,net647_c1,dummy48);
wire dummy49;
SPLITT SplitCLK_2_568(net944,net646_c1,dummy49);
wire dummy50;
SPLITT SplitCLK_2_569(net1176,net645_c1,dummy50);
wire dummy51;
SPLITT SplitCLK_2_570(net1138,net644_c1,dummy51);
wire dummy52;
SPLITT SplitCLK_2_571(net1075,net643_c1,dummy52);
wire dummy53;
SPLITT SplitCLK_2_572(net850,net642_c1,dummy53);
wire dummy54;
SPLITT SplitCLK_4_573(net838,net641_c1,dummy54);
wire dummy55;
SPLITT SplitCLK_4_574(net1108,net640_c1,dummy55);
wire dummy56;
SPLITT SplitCLK_2_575(net1064,net639_c1,dummy56);
wire dummy57;
SPLITT SplitCLK_4_576(net1171,net638_c1,dummy57);
wire dummy58;
SPLITT SplitCLK_2_577(net972,net637_c1,dummy58);
wire dummy59;
SPLITT SplitCLK_4_578(net1111,net636_c1,dummy59);
wire dummy60;
SPLITT SplitCLK_4_579(net998,net635_c1,dummy60);
wire dummy61;
SPLITT SplitCLK_2_580(net1010,net634_c1,dummy61);
wire dummy62;
SPLITT SplitCLK_2_581(net1060,net633_c1,dummy62);
wire dummy63;
SPLITT SplitCLK_2_582(net1072,net632_c1,dummy63);
wire dummy64;
SPLITT SplitCLK_4_583(net1061,net631_c1,dummy64);
wire dummy65;
SPLITT SplitCLK_4_584(net874,net630_c1,dummy65);
wire dummy66;
SPLITT SplitCLK_2_585(net942,net629_c1,dummy66);
wire dummy67;
SPLITT SplitCLK_4_586(net943,net628_c1,dummy67);
wire dummy68;
SPLITT SplitCLK_4_587(net918,net627_c1,dummy68);
wire dummy69;
SPLITT SplitCLK_4_588(net1114,net626_c1,dummy69);
wire dummy70;
SPLITT SplitCLK_4_589(net1028,net625_c1,dummy70);
wire dummy71;
SPLITT SplitCLK_4_590(net815,net624_c1,dummy71);
wire dummy72;
SPLITT SplitCLK_2_591(net1186,net623_c1,dummy72);
wire dummy73;
SPLITT SplitCLK_2_592(net746,net622_c1,dummy73);
wire dummy74;
SPLITT SplitCLK_4_593(net852,net621_c1,dummy74);
wire dummy75;
SPLITT SplitCLK_4_594(net1132,net620_c1,dummy75);
wire dummy76;
SPLITT SplitCLK_4_595(net1192,net619_c1,dummy76);
wire dummy77;
SPLITT SplitCLK_2_596(net882,net618_c1,dummy77);
wire dummy78;
SPLITT SplitCLK_4_597(net776,net617_c1,dummy78);
wire dummy79;
SPLITT SplitCLK_4_598(net987,net616_c1,dummy79);
wire dummy80;
SPLITT SplitCLK_2_599(net802,net615_c1,dummy80);
wire dummy81;
SPLITT SplitCLK_4_600(net1004,net614_c1,dummy81);
wire dummy82;
SPLITT SplitCLK_4_601(net899,net613_c1,dummy82);
wire dummy83;
SPLITT SplitCLK_4_602(net1002,net612_c1,dummy83);
wire dummy84;
SPLITT SplitCLK_4_603(net1016,net611_c1,dummy84);
wire dummy85;
SPLITT SplitCLK_4_604(net808,net610_c1,dummy85);
wire dummy86;
SPLITT SplitCLK_2_605(net816,net609_c1,dummy86);
wire dummy87;
SPLITT SplitCLK_2_606(net790,net608_c1,dummy87);
wire dummy88;
SPLITT SplitCLK_4_607(net752,net607_c1,dummy88);
wire dummy89;
SPLITT SplitCLK_2_608(net744,net606_c1,dummy89);
wire dummy90;
SPLITT SplitCLK_2_609(net806,net605_c1,dummy90);
wire dummy91;
SPLITT SplitCLK_4_610(net900,net604_c1,dummy91);
wire dummy92;
SPLITT SplitCLK_2_611(net809,net603_c1,dummy92);
wire dummy93;
SPLITT SplitCLK_2_612(net740,net602_c1,dummy93);
wire dummy94;
SPLITT SplitCLK_2_613(net784,net601_c1,dummy94);
wire dummy95;
SPLITT SplitCLK_4_614(net866,net600_c1,dummy95);
wire dummy96;
SPLITT SplitCLK_4_615(net772,net599_c1,dummy96);
wire dummy97;
SPLITT SplitCLK_4_616(net773,net598_c1,dummy97);
wire dummy98;
SPLITT SplitCLK_4_617(net1203,net597_c1,dummy98);
wire dummy99;
SPLITT SplitCLK_4_618(net842,net596_c1,dummy99);
wire dummy100;
SPLITT SplitCLK_2_619(net722,net595_c1,dummy100);
wire dummy101;
SPLITT SplitCLK_4_620(net770,net594_c1,dummy101);
wire dummy102;
SPLITT SplitCLK_2_621(net1003,net593_c1,dummy102);
wire dummy103;
SPLITT SplitCLK_2_622(net858,net592_c1,dummy103);
wire dummy104;
SPLITT SplitCLK_4_623(net741,net591_c1,dummy104);
wire dummy105;
SPLITT SplitCLK_2_624(net739,net590_c1,dummy105);
wire dummy106;
SPLITT SplitCLK_4_625(net724,net589_c1,dummy106);
wire dummy107;
SPLITT SplitCLK_4_626(net747,net588_c1,dummy107);
wire dummy108;
SPLITT SplitCLK_2_627(net820,net587_c1,dummy108);
wire dummy109;
SPLITT SplitCLK_2_628(net725,net586_c1,dummy109);
wire dummy110;
SPLITT SplitCLK_4_629(net928,net585_c1,dummy110);
wire dummy111;
SPLITT SplitCLK_4_630(net786,net584_c1,dummy111);
wire dummy112;
SPLITT SplitCLK_4_631(net1208,net583_c1,dummy112);
wire dummy113;
SPLITT SplitCLK_2_632(net915,net582_c1,dummy113);
wire dummy114;
SPLITT SplitCLK_4_633(net921,net581_c1,dummy114);
wire dummy115;
SPLITT SplitCLK_4_634(net982,net580_c1,dummy115);
wire dummy116;
SPLITT SplitCLK_2_635(net1017,net579_c1,dummy116);
wire dummy117;
SPLITT SplitCLK_4_636(net728,net578_c1,dummy117);
wire dummy118;
SPLITT SplitCLK_2_637(net929,net577_c1,dummy118);
wire dummy119;
SPLITT SplitCLK_2_638(net1177,net576_c1,dummy119);
wire dummy120;
SPLITT SplitCLK_4_639(net1164,net575_c1,dummy120);
wire dummy121;
SPLITT SplitCLK_2_640(net1201,net574_c1,dummy121);
wire dummy122;
SPLITT SplitCLK_4_641(net716,net573_c1,dummy122);
wire dummy123;
SPLITT SplitCLK_2_642(net800,net572_c1,dummy123);
wire dummy124;
SPLITT SplitCLK_4_643(net730,net571_c1,dummy124);
wire dummy125;
SPLITT SplitCLK_4_644(net883,net570_c1,dummy125);
wire dummy126;
SPLITT SplitCLK_4_645(net754,net569_c1,dummy126);
wire dummy127;
SPLITT SplitCLK_2_646(net745,net568_c1,dummy127);
wire dummy128;
SPLITT SplitCLK_4_647(net1195,net567_c1,dummy128);
wire dummy129;
SPLITT SplitCLK_2_648(net1139,net566_c1,dummy129);
wire dummy130;
SPLITT SplitCLK_4_649(net779,net565_c1,dummy130);
wire dummy131;
SPLITT SplitCLK_2_650(net729,net564_c1,dummy131);
wire dummy132;
SPLITT SplitCLK_4_651(net1097,net563_c1,dummy132);
wire dummy133;
SPLITT SplitCLK_2_652(net1005,net562_c1,dummy133);
wire dummy134;
SPLITT SplitCLK_4_653(net881,net561_c1,dummy134);
wire dummy135;
SPLITT SplitCLK_2_654(net1115,net560_c1,dummy135);
wire dummy136;
SPLITT SplitCLK_4_655(net1011,net559_c1,dummy136);
wire dummy137;
SPLITT SplitCLK_2_656(net973,net558_c1,dummy137);
wire dummy138;
SPLITT SplitCLK_2_657(net1018,net557_c1,dummy138);
wire dummy139;
SPLITT SplitCLK_2_658(net996,net556_c1,dummy139);
wire dummy140;
SPLITT SplitCLK_2_659(net803,net555_c1,dummy140);
wire dummy141;
SPLITT SplitCLK_4_660(net1065,net554_c1,dummy141);
wire dummy142;
SPLITT SplitCLK_2_661(net1059,net553_c1,dummy142);
wire dummy143;
SPLITT SplitCLK_4_662(net1012,net552_c1,dummy143);
wire dummy144;
SPLITT SplitCLK_2_663(net1188,net551_c1,dummy144);
wire dummy145;
SPLITT SplitCLK_4_664(net844,net550_c1,dummy145);
wire dummy146;
SPLITT SplitCLK_2_665(net1048,net549_c1,dummy146);
wire dummy147;
SPLITT SplitCLK_2_666(net1030,net548_c1,dummy147);
wire dummy148;
SPLITT SplitCLK_2_667(net731,net547_c1,dummy148);
wire dummy149;
SPLITT SplitCLK_4_668(net983,net546_c1,dummy149);
wire dummy150;
SPLITT SplitCLK_2_669(net851,net545_c1,dummy150);
wire dummy151;
SPLITT SplitCLK_4_670(net868,net544_c1,dummy151);
wire dummy152;
SPLITT SplitCLK_2_671(net807,net543_c1,dummy152);
wire dummy153;
SPLITT SplitCLK_2_672(net1078,net542_c1,dummy153);
wire dummy154;
SPLITT SplitCLK_4_673(net821,net541_c1,dummy154);
wire dummy155;
SPLITT SplitCLK_2_674(net867,net540_c1,dummy155);
wire dummy156;
SPLITT SplitCLK_4_675(net760,net539_c1,dummy156);
wire dummy157;
SPLITT SplitCLK_4_676(net1066,net538_c1,dummy157);
wire dummy158;
SPLITT SplitCLK_2_677(net753,net537_c1,dummy158);
wire dummy159;
SPLITT SplitCLK_4_678(net1019,net536_c1,dummy159);
wire dummy160;
SPLITT SplitCLK_2_679(net777,net535_c1,dummy160);
wire dummy161;
SPLITT SplitCLK_4_680(net801,net534_c1,dummy161);
wire dummy162;
SPLITT SplitCLK_2_681(net845,net533_c1,dummy162);
wire dummy163;
SPLITT SplitCLK_4_682(net873,net532_c1,dummy163);
wire dummy164;
SPLITT SplitCLK_4_683(net1049,net531_c1,dummy164);
wire dummy165;
SPLITT SplitCLK_2_684(net856,net530_c1,dummy165);
wire dummy166;
SPLITT SplitCLK_2_685(net836,net529_c1,dummy166);
wire dummy167;
SPLITT SplitCLK_4_686(net1031,net528_c1,dummy167);
wire dummy168;
SPLITT SplitCLK_2_687(net714,net527_c1,dummy168);
wire dummy169;
SPLITT SplitCLK_2_688(net980,net526_c1,dummy169);
wire dummy170;
SPLITT SplitCLK_4_689(net907,net525_c1,dummy170);
wire dummy171;
SPLITT SplitCLK_2_690(net869,net524_c1,dummy171);
wire dummy172;
SPLITT SplitCLK_2_691(net886,net523_c1,dummy172);
wire dummy173;
SPLITT SplitCLK_2_692(net1050,net522_c1,dummy173);
wire dummy174;
SPLITT SplitCLK_4_693(net1165,net521_c1,dummy174);
wire dummy175;
SPLITT SplitCLK_2_694(net857,net520_c1,dummy175);
wire dummy176;
SPLITT SplitCLK_2_695(net934,net519_c1,dummy176);
wire dummy177;
SPLITT SplitCLK_2_696(net1013,net518_c1,dummy177);
wire dummy178;
SPLITT SplitCLK_2_697(net1042,net517_c1,dummy178);
wire dummy179;
SPLITT SplitCLK_2_698(net717,net516_c1,dummy179);
wire dummy180;
SPLITT SplitCLK_4_699(net968,net515_c1,dummy180);
wire dummy181;
SPLITT SplitCLK_4_700(net1127,net514_c1,dummy181);
wire dummy182;
SPLITT SplitCLK_4_701(net887,net513_c1,dummy182);
wire dummy183;
SPLITT SplitCLK_2_702(net1095,net512_c1,dummy183);
wire dummy184;
SPLITT SplitCLK_4_703(net1051,net511_c1,dummy184);
wire dummy185;
SPLITT SplitCLK_4_704(net1189,net510_c1,dummy185);
wire dummy186;
SPLITT SplitCLK_4_705(net945,net509_c1,dummy186);
wire dummy187;
SPLITT SplitCLK_4_706(net1044,net508_c1,dummy187);
wire dummy188;
SPLITT SplitCLK_4_707(net761,net507_c1,dummy188);
wire dummy189;
SPLITT SplitCLK_4_708(net966,net506_c1,dummy189);
wire dummy190;
SPLITT SplitCLK_2_709(net1187,net505_c1,dummy190);
wire dummy191;
SPLITT SplitCLK_4_710(net1144,net504_c1,dummy191);
wire dummy192;
SPLITT SplitCLK_2_711(net875,net503_c1,dummy192);
wire dummy193;
SPLITT SplitCLK_2_712(net787,net502_c1,dummy193);
wire dummy194;
SPLITT SplitCLK_2_713(net1079,net501_c1,dummy194);
wire dummy195;
SPLITT SplitCLK_2_714(net1163,net500_c1,dummy195);
wire dummy196;
SPLITT SplitCLK_2_715(net919,net499_c1,dummy196);
wire dummy197;
SPLITT SplitCLK_2_716(net1206,net498_c1,dummy197);
wire dummy198;
SPLITT SplitCLK_4_717(net785,net497_c1,dummy198);
wire dummy199;
SPLITT SplitCLK_4_718(net1045,net496_c1,dummy199);
wire dummy200;
SPLITT SplitCLK_4_719(net759,net495_c1,dummy200);
wire dummy201;
SPLITT SplitCLK_4_720(net1207,net494_c1,dummy201);
wire dummy202;
SPLITT SplitCLK_2_721(net1146,net493_c1,dummy202);
wire dummy203;
SPLITT SplitCLK_4_722(net723,net492_c1,dummy203);
wire dummy204;
SPLITT SplitCLK_4_723(net791,net491_c1,dummy204);
wire dummy205;
SPLITT SplitCLK_4_724(net1178,net490_c1,dummy205);
wire dummy206;
SPLITT SplitCLK_4_725(net837,net489_c1,dummy206);
wire dummy207;
SPLITT SplitCLK_4_726(net1116,net488_c1,dummy207);
wire dummy208;
SPLITT SplitCLK_2_727(net1043,net487_c1,dummy208);
wire dummy209;
SPLITT SplitCLK_2_728(net853,net486_c1,dummy209);
wire dummy210;
SPLITT SplitCLK_4_729(net1147,net485_c1,dummy210);
wire dummy211;
SPLITT SplitCLK_4_730(net948,net484_c1,dummy211);
wire dummy212;
SPLITT SplitCLK_4_731(net710,net483_c1,dummy212);
wire dummy213;
SPLITT SplitCLK_2_732(net793,net482_c1,dummy213);
wire dummy214;
SPLITT SplitCLK_4_733(net859,net481_c1,dummy214);
wire dummy215;
SPLITT SplitCLK_4_734(net974,net480_c1,dummy215);
wire dummy216;
SPLITT SplitCLK_4_735(net1117,net479_c1,dummy216);
wire dummy217;
SPLITT SplitCLK_2_736(net1193,net478_c1,dummy217);
wire dummy218;
SPLITT SplitCLK_4_737(net950,net477_c1,dummy218);
wire dummy219;
SPLITT SplitCLK_2_738(net981,net476_c1,dummy219);
wire dummy220;
SPLITT SplitCLK_2_739(net711,net475_c1,dummy220);
wire dummy221;
SPLITT SplitCLK_4_740(net901,net474_c1,dummy221);
wire dummy222;
SPLITT SplitCLK_4_741(net997,net473_c1,dummy222);
wire dummy223;
SPLITT SplitCLK_2_742(net839,net472_c1,dummy223);
wire dummy224;
SPLITT SplitCLK_2_743(net1179,net471_c1,dummy224);
wire dummy225;
SPLITT SplitCLK_4_744(net771,net470_c1,dummy225);
wire dummy226;
SPLITT SplitCLK_2_745(net843,net469_c1,dummy226);
wire dummy227;
SPLITT SplitCLK_2_746(net1145,net468_c1,dummy227);
wire dummy228;
SPLITT SplitCLK_2_747(net1125,net467_c1,dummy228);
wire dummy229;
SPLITT SplitCLK_2_748(net975,net466_c1,dummy229);
wire dummy230;
SPLITT SplitCLK_4_749(net708,net465_c1,dummy230);
wire dummy231;
SPLITT SplitCLK_4_750(net1036,net464_c1,dummy231);
wire dummy232;
SPLITT SplitCLK_4_751(net817,net463_c1,dummy232);
wire dummy233;
SPLITT SplitCLK_2_752(net1133,net462_c1,dummy233);
wire dummy234;
SPLITT SplitCLK_4_753(net935,net461_c1,dummy234);
wire dummy235;
SPLITT SplitCLK_2_754(net1029,net460_c1,dummy235);
wire dummy236;
SPLITT SplitCLK_2_755(net709,net459_c1,dummy236);
wire dummy237;
SPLITT SplitCLK_4_756(net1037,net458_c1,dummy237);
wire dummy238;
SPLITT SplitCLK_2_757(net1109,net457_c1,dummy238);
wire dummy239;
SPLITT SplitCLK_4_758(net1131,net456_c1,dummy239);
wire dummy240;
SPLITT SplitCLK_2_759(net949,net455_c1,dummy240);
wire dummy241;
SPLITT SplitCLK_4_760(net989,net454_c1,dummy241);
wire dummy242;
SPLITT SplitCLK_4_761(net715,net453_c1,dummy242);
wire dummy243;
SPLITT SplitCLK_4_762(net1034,net452_c1,dummy243);
wire dummy244;
SPLITT SplitCLK_2_763(net1035,net451_c1,dummy244);
wire dummy245;
SPLITT SplitCLK_2_764(net999,net450_c1,dummy245);
wire dummy246;
SPLITT SplitCLK_4_765(net1073,net449_c1,dummy246);
wire dummy247;
SPLITT SplitCLK_4_766(net822,net448_c1,dummy247);
wire dummy248;
SPLITT SplitCLK_2_767(net967,net447_c1,dummy248);
wire dummy249;
SPLITT SplitCLK_4_768(net1067,net446_c1,dummy249);
wire dummy250;
SPLITT SplitCLK_2_769(net969,net445_c1,dummy250);
wire dummy251;
SPLITT SplitCLK_4_770(net755,net444_c1,dummy251);
SPLITT SplitCLK_0_771(net1212,net442_c1,net443_c1);
wire dummy252;
SPLITT Split_HOLD_869(net383,dummy252,net1213_c1);
wire dummy253;
SPLITT Split_HOLD_870(net426,dummy253,net1214_c1);
wire dummy254;
SPLITT Split_HOLD_871(net75,dummy254,net1215_c1);
wire dummy255;
SPLITT Split_HOLD_872(net306,dummy255,net1216_c1);
wire dummy256;
SPLITT Split_HOLD_873(net394,dummy256,net1217_c1);
wire dummy257;
SPLITT Split_HOLD_874(net408,dummy257,net1218_c1);
wire dummy258;
SPLITT Split_HOLD_875(net387,dummy258,net1219_c1);
wire dummy259;
SPLITT Split_HOLD_876(net420,dummy259,net1220_c1);
wire dummy260;
SPLITT Split_HOLD_877(net320,dummy260,net1221_c1);
INTERCONNECT TMS_Pad_Split_268_n727(TMS_Pad,net0);
INTERCONNECT NOTT_14_n50_AND2T_18_n54(net1_c1,net1);
INTERCONNECT AND2T_15_n51_Split_273_n732(net2_c1,net2);
INTERCONNECT NOTT_24_n60_Split_280_n739(net3_c1,net3);
INTERCONNECT NOTT_16_n52_DFFT_149__FPB_n608(net4_c1,net4);
INTERCONNECT AND2T_8_n44_DFFT_147__FPB_n606(net5_c1,net5);
INTERCONNECT NOTT_25_n61_Split_281_n740(net6_c1,net6);
INTERCONNECT AND2T_17_n53_OR2T_22_n58(net7_c1,net7);
INTERCONNECT NOTT_9_n45_AND2T_109_n151(net8_c1,net8);
INTERCONNECT OR2T_34_n70_Split_294_n753(net9_c1,net9);
INTERCONNECT NOTT_26_n62_Split_284_n743(net10_c1,net10);
INTERCONNECT AND2T_18_n54_AND2T_17_n53(net11_c1,net11);
INTERCONNECT NOTT_10_n46_OR2T_11_n47(net12_c1,net12);
INTERCONNECT AND2T_35_n71_DFFT_179__FPB_n638(net13_c1,net13);
INTERCONNECT AND2T_27_n63_Split_286_n745(net14_c1,net14);
INTERCONNECT AND2T_19_n55_Split_274_n733(net15_c1,net15);
INTERCONNECT OR2T_11_n47_DFFT_132__FPB_n591(net16_c1,net16);
INTERCONNECT AND2T_44_n80_Split_301_n760(net17_c1,net17);
INTERCONNECT AND2T_36_n72_Split_295_n754(net18_c1,net18);
INTERCONNECT AND2T_28_n64_DFFT_159__FPB_n618(net19_c1,net19);
INTERCONNECT AND2T_20_n56_Split_275_n734(net20_c1,net20);
INTERCONNECT NOTT_12_n48_Split_270_n729(net21_c1,net21);
INTERCONNECT OR2T_45_n81_OR2T_46_n82(net22_c1,net22);
INTERCONNECT AND2T_37_n73_OR2T_40_n76(net23_c1,net23);
INTERCONNECT AND2T_29_n65_Split_289_n748(net24_c1,net24);
INTERCONNECT OR2T_21_n57_DFFT_155__FPB_n614(net25_c1,net25);
INTERCONNECT AND2T_13_n49_AND2T_53_n89(net26_c1,net26);
INTERCONNECT OR2T_54_n90_AND2T_55_n91(net27_c1,net27);
INTERCONNECT OR2T_46_n82_OR2T_47_n83(net28_c1,net28);
INTERCONNECT AND2T_38_n74_AND2T_39_n75(net29_c1,net29);
INTERCONNECT AND2T_30_n66_DFFT_158__FPB_n617(net30_c1,net30);
INTERCONNECT OR2T_22_n58_DFFT_138__FPB_n597(net31_c1,net31);
INTERCONNECT AND2T_55_n91_OR2T_56_n92(net32_c1,net32);
INTERCONNECT OR2T_47_n83_OR2T_57_n93(net33_c1,net33);
INTERCONNECT AND2T_39_n75_OR2T_40_n76(net34_c1,net34);
INTERCONNECT AND2T_31_n67_Split_291_n750(net35_c1,net35);
INTERCONNECT NOTT_23_n59_Split_277_n736(net36_c1,net36);
INTERCONNECT OR2T_56_n92_OR2T_57_n93(net37_c1,net37);
INTERCONNECT AND2T_48_n84_OR2T_50_n86(net38_c1,net38);
INTERCONNECT OR2T_40_n76_Split_297_n756(net39_c1,net39);
INTERCONNECT AND2T_32_n68_OR2T_33_n69(net40_c1,net40);
INTERCONNECT OR2T_57_n93_OR2T_58_n94(net41_c1,net41);
INTERCONNECT AND2T_49_n85_OR2T_50_n86(net42_c1,net42);
INTERCONNECT AND2T_41_n77_Split_298_n757(net43_c1,net43);
INTERCONNECT OR2T_33_n69_OR2T_34_n70(net44_c1,net44);
INTERCONNECT OR2T_58_n94_AND2T_59_n95(net45_c1,net45);
INTERCONNECT OR2T_50_n86_Split_302_n761(net46_c1,net46);
INTERCONNECT AND2T_42_n78_OR2T_46_n82(net47_c1,net47);
INTERCONNECT AND2T_59_n95_DFFT_123__FBL_n582(net48_c1,net48);
INTERCONNECT AND2T_51_n87_OR2T_56_n92(net49_c1,net49);
INTERCONNECT AND2T_43_n79_Split_300_n759(net50_c1,net50);
INTERCONNECT OR2T_60_n96_Split_304_n763(net51_c1,net51);
INTERCONNECT AND2T_52_n88_Split_303_n762(net52_c1,net52);
INTERCONNECT OR2T_61_n97_AND2T_62_n98(net53_c1,net53);
INTERCONNECT AND2T_53_n89_OR2T_54_n90(net54_c1,net54);
INTERCONNECT AND2T_62_n98_OR2T_71_n107(net55_c1,net55);
INTERCONNECT AND2T_63_n99_OR2T_64_n100(net56_c1,net56);
INTERCONNECT OR2T_64_n100_Split_305_n764(net57_c1,net57);
INTERCONNECT AND2T_65_n101_DFFT_199__FPB_n658(net58_c1,net58);
INTERCONNECT AND2T_74_n110_Split_309_n768(net59_c1,net59);
INTERCONNECT AND2T_66_n102_Split_306_n765(net60_c1,net60);
INTERCONNECT XOR2T_75_n111_DFFT_209__FPB_n668(net61_c1,net61);
INTERCONNECT AND2T_67_n103_Split_307_n766(net62_c1,net62);
INTERCONNECT OR2T_84_n120_OR2T_88_n124(net63_c1,net63);
INTERCONNECT AND2T_76_n112_DFFT_212__FPB_n671(net64_c1,net64);
INTERCONNECT OR2T_68_n104_OR2T_69_n105(net65_c1,net65);
INTERCONNECT AND2T_85_n121_AND2T_86_n122(net66_c1,net66);
INTERCONNECT AND2T_77_n113_Split_310_n769(net67_c1,net67);
INTERCONNECT OR2T_69_n105_OR2T_70_n106(net68_c1,net68);
INTERCONNECT AND2T_94_n130_OR2T_96_n132(net69_c1,net69);
INTERCONNECT AND2T_86_n122_DFFT_215__FPB_n674(net70_c1,net70);
INTERCONNECT AND2T_78_n114_OR2T_79_n115(net71_c1,net71);
INTERCONNECT OR2T_70_n106_OR2T_71_n107(net72_c1,net72);
INTERCONNECT OR2T_95_n131_AND2T_94_n130(net73_c1,net73);
INTERCONNECT OR2T_87_n123_OR2T_88_n124(net74_c1,net74);
INTERCONNECT OR2T_79_n115_Split_HOLD_871(net75_c1,net75);
INTERCONNECT OR2T_71_n107_AND2T_72_n108(net76_c1,net76);
INTERCONNECT OR2T_96_n132_OR2T_97_n133(net77_c1,net77);
INTERCONNECT OR2T_88_n124_OR2T_89_n125(net78_c1,net78);
INTERCONNECT OR2T_80_n116_OR2T_89_n125(net79_c1,net79);
INTERCONNECT AND2T_72_n108_Split_308_n767(net80_c1,net80);
INTERCONNECT OR2T_97_n133_OR2T_98_n134(net81_c1,net81);
INTERCONNECT OR2T_89_n125_AND2T_90_n126(net82_c1,net82);
INTERCONNECT AND2T_81_n117_AND2T_82_n118(net83_c1,net83);
INTERCONNECT AND2T_73_n109_DFFT_213__FPB_n672(net84_c1,net84);
INTERCONNECT AND2T_108_n150_Split_318_n777(net85_c1,net85);
INTERCONNECT OR2T_98_n134_OR2T_99_n135(net86_c1,net86);
INTERCONNECT AND2T_90_n126_Split_311_n770(net87_c1,net87);
INTERCONNECT AND2T_82_n118_OR2T_83_n119(net88_c1,net88);
INTERCONNECT AND2T_109_n151_Split_321_n780(net89_c1,net89);
INTERCONNECT OR2T_99_n135_AND2T_100_n136(net90_c1,net90);
INTERCONNECT AND2T_91_n127_DFFT_231__FPB_n690(net91_c1,net91);
INTERCONNECT OR2T_83_n119_OR2T_84_n120(net92_c1,net92);
INTERCONNECT NOTT_112_n160_Split_330_n789(net93_c1,net93);
INTERCONNECT AND2T_110_n152_Split_324_n783(net94_c1,net94);
INTERCONNECT AND2T_100_n136_Split_314_n773(net95_c1,net95);
INTERCONNECT AND2T_92_n128_DFFT_230__FPB_n689(net96_c1,net96);
INTERCONNECT NOTT_111_n153_Split_327_n786(net97_c1,net97);
INTERCONNECT AND2T_93_n129_OR2T_96_n132(net98_c1,net98);
INTERCONNECT AND2T_107_n149_Split_315_n774(net99_c1,net99);
INTERCONNECT Split_341_n800_Split_343_n802(net100_c1,net100);
INTERCONNECT Split_342_n801_AND2T_29_n65(net101_c1,net101);
INTERCONNECT Split_351_n810_DFFT_238__FPB_n697(net102_c1,net102);
INTERCONNECT Split_343_n802_DFFT_157__FPB_n616(net103_c1,net103);
INTERCONNECT Split_271_n730_AND2T_15_n51(net104_c1,net104);
INTERCONNECT TRST_Pad_NOTT_23_n59(TRST_Pad,net105);
INTERCONNECT Split_352_n811_Split_354_n813(net106_c1,net106);
INTERCONNECT Split_344_n803_Split_346_n805(net107_c1,net107);
INTERCONNECT Split_272_n731_AND2T_108_n150(net108_c1,net108);
INTERCONNECT Split_281_n740_Split_283_n742(net109_c1,net109);
INTERCONNECT Split_345_n804_DFFT_208__FPB_n667(net110_c1,net110);
INTERCONNECT Split_273_n732_DFFT_207__FPB_n666(net111_c1,net111);
INTERCONNECT Split_353_n812_AND2T_20_n56(net112_c1,net112);
INTERCONNECT Split_346_n805_DFFT_227__FPB_n686(net113_c1,net113);
INTERCONNECT Split_274_n733_AND2T_93_n129(net114_c1,net114);
INTERCONNECT Split_354_n813_DFFT_153__FPB_n612(net115_c1,net115);
INTERCONNECT Split_282_n741_AND2T_36_n72(net116_c1,net116);
INTERCONNECT Split_355_n814_Split_357_n816(net117_c1,net117);
INTERCONNECT Split_291_n750_Split_293_n752(net118_c1,net118);
INTERCONNECT Split_275_n734_Split_276_n735(net119_c1,net119);
INTERCONNECT Split_347_n806_DFFT_239__FPB_n698(net120_c1,net120);
INTERCONNECT Split_283_n742_OR2T_95_n131(net121_c1,net121);
INTERCONNECT Split_348_n807_Split_350_n809(net122_c1,net122);
INTERCONNECT Split_268_n727_Split_269_n728(net123_c1,net123);
INTERCONNECT Split_284_n743_Split_285_n744(net124_c1,net124);
INTERCONNECT Split_276_n735_DFFT_175__FPB_n634(net125_c1,net125);
INTERCONNECT Split_292_n751_AND2T_52_n88(net126_c1,net126);
INTERCONNECT Split_356_n815_NOTT_9_n45(net127_c1,net127);
INTERCONNECT Split_277_n736_Split_279_n738(net128_c1,net128);
INTERCONNECT Split_269_n728_DFFT_113__FPB_n164(net129_c1,net129);
INTERCONNECT Split_293_n752_AND2T_66_n102(net130_c1,net130);
INTERCONNECT Split_301_n760_OR2T_64_n100(net131_c1,net131);
INTERCONNECT Split_285_n744_AND2T_31_n67(net132_c1,net132);
INTERCONNECT Split_349_n808_AND2T_29_n65(net133_c1,net133);
INTERCONNECT Split_357_n816_DFFT_148__FPB_n607(net134_c1,net134);
INTERCONNECT Split_286_n745_Split_288_n747(net135_c1,net135);
INTERCONNECT Split_270_n729_Split_272_n731(net136_c1,net136);
INTERCONNECT Split_278_n737_DFFT_200__FPB_n659(net137_c1,net137);
INTERCONNECT Split_350_n809_DFFT_166__FPB_n625(net138_c1,net138);
INTERCONNECT Split_302_n761_OR2T_84_n120(net139_c1,net139);
INTERCONNECT Split_294_n753_OR2T_61_n97(net140_c1,net140);
INTERCONNECT Split_311_n770_Split_313_n772(net141_c1,net141);
INTERCONNECT Split_279_n738_DFFT_232__FPB_n691(net142_c1,net142);
INTERCONNECT Split_303_n762_OR2T_60_n96(net143_c1,net143);
INTERCONNECT Split_295_n754_Split_296_n755(net144_c1,net144);
INTERCONNECT Split_287_n746_AND2T_43_n79(net145_c1,net145);
INTERCONNECT Split_312_n771_DFFT_143__FPB_n602(net146_c1,net146);
INTERCONNECT Split_304_n763_DFFT_187__FPB_n646(net147_c1,net147);
INTERCONNECT Split_280_n739_DFFT_211__FPB_n670(net148_c1,net148);
INTERCONNECT Split_288_n747_AND2T_53_n89(net149_c1,net149);
INTERCONNECT Split_296_n755_AND2T_41_n77(net150_c1,net150);
INTERCONNECT Split_321_n780_Split_323_n782(net151_c1,net151);
INTERCONNECT Split_289_n748_Split_290_n749(net152_c1,net152);
INTERCONNECT Split_313_n772_DFFT_146__FPB_n605(net153_c1,net153);
INTERCONNECT Split_297_n756_DFFT_170__FPB_n629(net154_c1,net154);
INTERCONNECT Split_305_n764_AND2T_91_n127(net155_c1,net155);
INTERCONNECT Split_298_n757_Split_299_n758(net156_c1,net156);
INTERCONNECT Split_314_n773_DFFT_145__FPB_n604(net157_c1,net157);
INTERCONNECT Split_306_n765_AND2T_73_n109(net158_c1,net158);
INTERCONNECT Split_290_n749_DFFT_171__FPB_n630(net159_c1,net159);
INTERCONNECT Split_322_n781_AND2T_28_n64(net160_c1,net160);
INTERCONNECT Split_315_n774_Split_317_n776(net161_c1,net161);
INTERCONNECT Split_307_n766_DFFT_198__FPB_n657(net162_c1,net162);
INTERCONNECT Split_299_n758_OR2T_83_n119(net163_c1,net163);
INTERCONNECT Split_323_n782_DFFT_196__FPB_n655(net164_c1,net164);
INTERCONNECT Split_331_n790_AND2T_13_n49(net165_c1,net165);
INTERCONNECT Split_324_n783_Split_326_n785(net166_c1,net166);
INTERCONNECT Split_308_n767_DFFT_127__FBL_n586(net167_c1,net167);
INTERCONNECT Split_300_n759_OR2T_60_n96(net168_c1,net168);
INTERCONNECT Split_332_n791_AND2T_107_n149(net169_c1,net169);
INTERCONNECT Split_316_n775_AND2T_32_n68(net170_c1,net170);
INTERCONNECT Split_333_n792_Split_335_n794(net171_c1,net171);
INTERCONNECT Split_309_n768_AND2T_86_n122(net172_c1,net172);
INTERCONNECT Split_317_n776_AND2T_49_n85(net173_c1,net173);
INTERCONNECT Split_325_n784_DFFT_154__FPB_n613(net174_c1,net174);
INTERCONNECT Split_318_n777_Split_320_n779(net175_c1,net175);
INTERCONNECT Split_326_n785_DFFT_169__FPB_n628(net176_c1,net176);
INTERCONNECT Split_310_n769_AND2T_92_n128(net177_c1,net177);
INTERCONNECT Split_334_n793_DFFT_167__FPB_n626(net178_c1,net178);
INTERCONNECT Split_327_n786_Split_329_n788(net179_c1,net179);
INTERCONNECT Split_335_n794_DFFT_188__FPB_n647(net180_c1,net180);
INTERCONNECT Split_319_n778_AND2T_41_n77(net181_c1,net181);
INTERCONNECT Split_336_n795_Split_338_n797(net182_c1,net182);
INTERCONNECT Split_320_n779_AND2T_63_n99(net183_c1,net183);
INTERCONNECT Split_328_n787_DFFT_160__FPB_n619(net184_c1,net184);
INTERCONNECT Split_329_n788_DFFT_193__FPB_n652(net185_c1,net185);
INTERCONNECT Split_337_n796_AND2T_85_n121(net186_c1,net186);
INTERCONNECT Split_330_n789_Split_332_n791(net187_c1,net187);
INTERCONNECT Split_338_n797_DFFT_225__FPB_n684(net188_c1,net188);
INTERCONNECT Split_339_n798_DFFT_103_state_obs2_buf(net189_c1,net189);
INTERCONNECT Split_340_n799_DFFT_150__FPB_n609(net190_c1,net190);
INTERCONNECT Split_341_n800_Split_342_n801(net191_c1,net191);
INTERCONNECT Split_342_n801_NOTT_25_n61(net192_c1,net192);
INTERCONNECT Split_271_n730_AND2T_13_n49(net193_c1,net193);
INTERCONNECT Split_343_n802_DFFT_105_state0_buf(net194_c1,net194);
INTERCONNECT Split_351_n810_AND2T_110_n152(net195_c1,net195);
INTERCONNECT Split_272_n731_AND2T_107_n149(net196_c1,net196);
INTERCONNECT Split_344_n803_Split_345_n804(net197_c1,net197);
INTERCONNECT Split_352_n811_Split_353_n812(net198_c1,net198);
INTERCONNECT Split_273_n732_AND2T_77_n113(net199_c1,net199);
INTERCONNECT Split_281_n740_Split_282_n741(net200_c1,net200);
INTERCONNECT Split_345_n804_DFFT_106_state1_buf(net201_c1,net201);
INTERCONNECT Split_353_n812_NOTT_12_n48(net202_c1,net202);
INTERCONNECT Split_274_n733_AND2T_82_n118(net203_c1,net203);
INTERCONNECT Split_282_n741_AND2T_27_n63(net204_c1,net204);
INTERCONNECT Split_346_n805_DFFT_214__FPB_n673(net205_c1,net205);
INTERCONNECT Split_354_n813_XOR2T_75_n111(net206_c1,net206);
INTERCONNECT Split_275_n734_DFFT_229__FPB_n688(net207_c1,net207);
INTERCONNECT Split_283_n742_AND2T_85_n121(net208_c1,net208);
INTERCONNECT Split_291_n750_Split_292_n751(net209_c1,net209);
INTERCONNECT Split_347_n806_AND2T_110_n152(net210_c1,net210);
INTERCONNECT Split_355_n814_Split_356_n815(net211_c1,net211);
INTERCONNECT Split_268_n727_DFFT_114__FPB_n165(net212_c1,net212);
INTERCONNECT Split_276_n735_AND2T_74_n110(net213_c1,net213);
INTERCONNECT Split_284_n743_OR2T_95_n131(net214_c1,net214);
INTERCONNECT Split_292_n751_AND2T_32_n68(net215_c1,net215);
INTERCONNECT Split_348_n807_Split_349_n808(net216_c1,net216);
INTERCONNECT Split_356_n815_AND2T_8_n44(net217_c1,net217);
INTERCONNECT Split_269_n728_NOTT_111_n153(net218_c1,net218);
INTERCONNECT Split_277_n736_Split_278_n737(net219_c1,net219);
INTERCONNECT Split_285_n744_AND2T_27_n63(net220_c1,net220);
INTERCONNECT Split_293_n752_AND2T_63_n99(net221_c1,net221);
INTERCONNECT Split_349_n808_NOTT_26_n62(net222_c1,net222);
INTERCONNECT Split_357_n816_AND2T_20_n56(net223_c1,net223);
INTERCONNECT Split_301_n760_OR2T_45_n81(net224_c1,net224);
INTERCONNECT Split_278_n737_DFFT_180__FPB_n639(net225_c1,net225);
INTERCONNECT Split_286_n745_Split_287_n746(net226_c1,net226);
INTERCONNECT Split_294_n753_AND2T_35_n71(net227_c1,net227);
INTERCONNECT Split_270_n729_Split_271_n730(net228_c1,net228);
INTERCONNECT Split_350_n809_DFFT_164__FPB_n623(net229_c1,net229);
INTERCONNECT Split_302_n761_AND2T_51_n87(net230_c1,net230);
INTERCONNECT Split_279_n738_DFFT_216__FPB_n675(net231_c1,net231);
INTERCONNECT Split_287_n746_AND2T_28_n64(net232_c1,net232);
INTERCONNECT Split_295_n754_AND2T_44_n80(net233_c1,net233);
INTERCONNECT Split_303_n762_OR2T_54_n90(net234_c1,net234);
INTERCONNECT Split_311_n770_Split_312_n771(net235_c1,net235);
INTERCONNECT Split_288_n747_AND2T_48_n84(net236_c1,net236);
INTERCONNECT Split_296_n755_AND2T_37_n73(net237_c1,net237);
INTERCONNECT Split_280_n739_AND2T_66_n102(net238_c1,net238);
INTERCONNECT Split_304_n763_OR2T_87_n123(net239_c1,net239);
INTERCONNECT Split_312_n771_DFFT_141__FPB_n600(net240_c1,net240);
INTERCONNECT Split_289_n748_DFFT_210__FPB_n669(net241_c1,net241);
INTERCONNECT Split_297_n756_OR2T_68_n104(net242_c1,net242);
INTERCONNECT Split_305_n764_AND2T_65_n101(net243_c1,net243);
INTERCONNECT Split_313_n772_DFFT_144__FPB_n603(net244_c1,net244);
INTERCONNECT Split_321_n780_Split_322_n781(net245_c1,net245);
INTERCONNECT Split_298_n757_DFFT_197__FPB_n656(net246_c1,net246);
INTERCONNECT Split_290_n749_AND2T_30_n66(net247_c1,net247);
INTERCONNECT Split_306_n765_AND2T_67_n103(net248_c1,net248);
INTERCONNECT Split_314_n773_DFFT_142__FPB_n601(net249_c1,net249);
INTERCONNECT Split_322_n781_OR2T_21_n57(net250_c1,net250);
INTERCONNECT Split_299_n758_AND2T_42_n78(net251_c1,net251);
INTERCONNECT Split_307_n766_OR2T_97_n133(net252_c1,net252);
INTERCONNECT Split_315_n774_Split_316_n775(net253_c1,net253);
INTERCONNECT Split_323_n782_AND2T_39_n75(net254_c1,net254);
INTERCONNECT Split_331_n790_NOTT_10_n46(net255_c1,net255);
INTERCONNECT Split_308_n767_DFFT_124__FBL_n583(net256_c1,net256);
INTERCONNECT Split_316_n775_NOTT_14_n50(net257_c1,net257);
INTERCONNECT Split_324_n783_Split_325_n784(net258_c1,net258);
INTERCONNECT Split_332_n791_AND2T_19_n55(net259_c1,net259);
INTERCONNECT Split_300_n759_OR2T_45_n81(net260_c1,net260);
INTERCONNECT Split_309_n768_AND2T_76_n112(net261_c1,net261);
INTERCONNECT Split_317_n776_AND2T_44_n80(net262_c1,net262);
INTERCONNECT Split_325_n784_AND2T_30_n66(net263_c1,net263);
INTERCONNECT Split_333_n792_Split_334_n793(net264_c1,net264);
INTERCONNECT Split_318_n777_Split_319_n778(net265_c1,net265);
INTERCONNECT Split_326_n785_DFFT_165__FPB_n624(net266_c1,net266);
INTERCONNECT Split_334_n793_NOTT_24_n60(net267_c1,net267);
INTERCONNECT Split_310_n769_AND2T_78_n114(net268_c1,net268);
INTERCONNECT Split_319_n778_NOTT_16_n52(net269_c1,net269);
INTERCONNECT Split_327_n786_Split_328_n787(net270_c1,net270);
INTERCONNECT Split_335_n794_DFFT_172__FPB_n631(net271_c1,net271);
INTERCONNECT Split_328_n787_AND2T_38_n74(net272_c1,net272);
INTERCONNECT Split_336_n795_Split_337_n796(net273_c1,net273);
INTERCONNECT Split_320_n779_AND2T_48_n84(net274_c1,net274);
INTERCONNECT Split_329_n788_DFFT_176__FPB_n635(net275_c1,net275);
INTERCONNECT Split_337_n796_AND2T_81_n117(net276_c1,net276);
INTERCONNECT Split_338_n797_DFFT_222__FPB_n681(net277_c1,net277);
INTERCONNECT Split_330_n789_Split_331_n790(net278_c1,net278);
INTERCONNECT Split_339_n798_AND2T_8_n44(net279_c1,net279);
INTERCONNECT Split_340_n799_DFFT_104_state_obs3_buf(net280_c1,net280);
INTERCONNECT DFFT_101_state_obs0_buf_DFFT_115__PIPL_n166(net281_c1,net281);
INTERCONNECT DFFT_102_state_obs1_buf_DFFT_116__PIPL_n167(net282_c1,net282);
INTERCONNECT DFFT_103_state_obs2_buf_DFFT_117__PIPL_n168(net283_c1,net283);
INTERCONNECT DFFT_104_state_obs3_buf_DFFT_118__PIPL_n169(net284_c1,net284);
INTERCONNECT DFFT_119__PIPL_n170_DFFT_101_state_obs0_buf(net285_c1,net285);
INTERCONNECT DFFT_120__PIPL_n171_DFFT_102_state_obs1_buf(net286_c1,net286);
INTERCONNECT DFFT_115__PIPL_n166_DFFT_240__FPB_n699(net287_c1,net287);
INTERCONNECT DFFT_116__PIPL_n167_DFFT_246__FPB_n705(net288_c1,net288);
INTERCONNECT DFFT_117__PIPL_n168_DFFT_252__FPB_n711(net289_c1,net289);
INTERCONNECT DFFT_118__PIPL_n169_DFFT_260__FPB_n719(net290_c1,net290);
INTERCONNECT DFFT_121__FBL_n580_Split_339_n798(net291_c1,net291);
INTERCONNECT DFFT_122__FBL_n581_Split_340_n799(net292_c1,net292);
INTERCONNECT DFFT_131__FBL_n590_Split_355_n814(net293_c1,net293);
INTERCONNECT DFFT_123__FBL_n582_Split_341_n800(net294_c1,net294);
INTERCONNECT DFFT_124__FBL_n583_Split_344_n803(net295_c1,net295);
INTERCONNECT DFFT_125__FBL_n584_XOR2T_75_n111(net296_c1,net296);
INTERCONNECT DFFT_126__FBL_n585_Split_347_n806(net297_c1,net297);
INTERCONNECT DFFT_127__FBL_n586_Split_348_n807(net298_c1,net298);
INTERCONNECT DFFT_128__FBL_n587_Split_351_n810(net299_c1,net299);
INTERCONNECT DFFT_129__FBL_n588_NOTT_112_n160(net300_c1,net300);
INTERCONNECT DFFT_130__FBL_n589_Split_352_n811(net301_c1,net301);
INTERCONNECT DFFT_113__FPB_n164_Split_333_n792(net302_c1,net302);
INTERCONNECT DFFT_114__FPB_n165_Split_336_n795(net303_c1,net303);
INTERCONNECT DFFT_141__FPB_n600_DFFT_125__FBL_n584(net304_c1,net304);
INTERCONNECT DFFT_142__FPB_n601_DFFT_126__FBL_n585(net305_c1,net305);
INTERCONNECT DFFT_151__FPB_n610_Split_HOLD_872(net306_c1,net306);
INTERCONNECT DFFT_143__FPB_n602_DFFT_128__FBL_n587(net307_c1,net307);
INTERCONNECT DFFT_144__FPB_n603_DFFT_129__FBL_n588(net308_c1,net308);
INTERCONNECT DFFT_152__FPB_n611_AND2T_18_n54(net309_c1,net309);
INTERCONNECT DFFT_241__FPB_n700_DFFT_242__FPB_n701(net310_c1,net310);
INTERCONNECT DFFT_161__FPB_n620_DFFT_162__FPB_n621(net311_c1,net311);
INTERCONNECT DFFT_145__FPB_n604_DFFT_130__FBL_n589(net312_c1,net312);
INTERCONNECT DFFT_153__FPB_n612_AND2T_19_n55(net313_c1,net313);
INTERCONNECT DFFT_242__FPB_n701_DFFT_243__FPB_n702(net314_c1,net314);
INTERCONNECT DFFT_162__FPB_n621_DFFT_163__FPB_n622(net315_c1,net315);
INTERCONNECT DFFT_146__FPB_n605_DFFT_131__FBL_n590(net316_c1,net316);
INTERCONNECT DFFT_154__FPB_n613_OR2T_21_n57(net317_c1,net317);
INTERCONNECT DFFT_243__FPB_n702_DFFT_244__FPB_n703(net318_c1,net318);
INTERCONNECT DFFT_155__FPB_n614_DFFT_156__FPB_n615(net319_c1,net319);
INTERCONNECT DFFT_171__FPB_n630_Split_HOLD_877(net320_c1,net320);
INTERCONNECT DFFT_163__FPB_n622_AND2T_35_n71(net321_c1,net321);
INTERCONNECT DFFT_147__FPB_n606_OR2T_11_n47(net322_c1,net322);
INTERCONNECT DFFT_252__FPB_n711_DFFT_253__FPB_n712(net323_c1,net323);
INTERCONNECT DFFT_244__FPB_n703_DFFT_245_state_obs0(net324_c1,net324);
INTERCONNECT DFFT_172__FPB_n631_DFFT_173__FPB_n632(net325_c1,net325);
INTERCONNECT DFFT_164__FPB_n623_AND2T_36_n72(net326_c1,net326);
INTERCONNECT DFFT_156__FPB_n615_OR2T_22_n58(net327_c1,net327);
INTERCONNECT DFFT_148__FPB_n607_AND2T_15_n51(net328_c1,net328);
INTERCONNECT DFFT_261__FPB_n720_DFFT_262__FPB_n721(net329_c1,net329);
INTERCONNECT DFFT_253__FPB_n712_DFFT_254__FPB_n713(net330_c1,net330);
INTERCONNECT DFFT_181__FPB_n640_DFFT_182__FPB_n641(net331_c1,net331);
INTERCONNECT DFFT_173__FPB_n632_DFFT_174__FPB_n633(net332_c1,net332);
INTERCONNECT DFFT_165__FPB_n624_AND2T_37_n73(net333_c1,net333);
INTERCONNECT DFFT_157__FPB_n616_AND2T_31_n67(net334_c1,net334);
INTERCONNECT DFFT_149__FPB_n608_AND2T_17_n53(net335_c1,net335);
INTERCONNECT DFFT_262__FPB_n721_DFFT_263__FPB_n722(net336_c1,net336);
INTERCONNECT DFFT_254__FPB_n713_DFFT_255__FPB_n714(net337_c1,net337);
INTERCONNECT DFFT_246__FPB_n705_DFFT_247__FPB_n706(net338_c1,net338);
INTERCONNECT DFFT_182__FPB_n641_DFFT_183__FPB_n642(net339_c1,net339);
INTERCONNECT DFFT_150__FPB_n609_DFFT_151__FPB_n610(net340_c1,net340);
INTERCONNECT DFFT_174__FPB_n633_AND2T_51_n87(net341_c1,net341);
INTERCONNECT DFFT_166__FPB_n625_AND2T_38_n74(net342_c1,net342);
INTERCONNECT DFFT_158__FPB_n617_OR2T_33_n69(net343_c1,net343);
INTERCONNECT DFFT_263__FPB_n722_DFFT_264__FPB_n723(net344_c1,net344);
INTERCONNECT DFFT_255__FPB_n714_DFFT_256__FPB_n715(net345_c1,net345);
INTERCONNECT DFFT_247__FPB_n706_DFFT_248__FPB_n707(net346_c1,net346);
INTERCONNECT DFFT_191__FPB_n650_DFFT_192__FPB_n651(net347_c1,net347);
INTERCONNECT DFFT_183__FPB_n642_DFFT_184__FPB_n643(net348_c1,net348);
INTERCONNECT DFFT_167__FPB_n626_DFFT_168__FPB_n627(net349_c1,net349);
INTERCONNECT DFFT_175__FPB_n634_AND2T_52_n88(net350_c1,net350);
INTERCONNECT DFFT_159__FPB_n618_OR2T_34_n70(net351_c1,net351);
INTERCONNECT DFFT_264__FPB_n723_DFFT_265__FPB_n724(net352_c1,net352);
INTERCONNECT DFFT_256__FPB_n715_DFFT_257__FPB_n716(net353_c1,net353);
INTERCONNECT DFFT_248__FPB_n707_DFFT_249__FPB_n708(net354_c1,net354);
INTERCONNECT DFFT_184__FPB_n643_DFFT_185__FPB_n644(net355_c1,net355);
INTERCONNECT DFFT_176__FPB_n635_DFFT_177__FPB_n636(net356_c1,net356);
INTERCONNECT DFFT_160__FPB_n619_DFFT_161__FPB_n620(net357_c1,net357);
INTERCONNECT DFFT_192__FPB_n651_AND2T_62_n98(net358_c1,net358);
INTERCONNECT DFFT_168__FPB_n627_AND2T_42_n78(net359_c1,net359);
INTERCONNECT DFFT_265__FPB_n724_DFFT_266__FPB_n725(net360_c1,net360);
INTERCONNECT DFFT_257__FPB_n716_DFFT_258__FPB_n717(net361_c1,net361);
INTERCONNECT DFFT_249__FPB_n708_DFFT_250__FPB_n709(net362_c1,net362);
INTERCONNECT DFFT_201__FPB_n660_DFFT_202__FPB_n661(net363_c1,net363);
INTERCONNECT DFFT_193__FPB_n652_DFFT_194__FPB_n653(net364_c1,net364);
INTERCONNECT DFFT_185__FPB_n644_DFFT_186__FPB_n645(net365_c1,net365);
INTERCONNECT DFFT_177__FPB_n636_DFFT_178__FPB_n637(net366_c1,net366);
INTERCONNECT DFFT_169__FPB_n628_AND2T_43_n79(net367_c1,net367);
INTERCONNECT DFFT_266__FPB_n725_DFFT_267_state_obs3(net368_c1,net368);
INTERCONNECT DFFT_258__FPB_n717_DFFT_259_state_obs2(net369_c1,net369);
INTERCONNECT DFFT_250__FPB_n709_DFFT_251_state_obs1(net370_c1,net370);
INTERCONNECT DFFT_202__FPB_n661_DFFT_203__FPB_n662(net371_c1,net371);
INTERCONNECT DFFT_194__FPB_n653_DFFT_195__FPB_n654(net372_c1,net372);
INTERCONNECT DFFT_186__FPB_n645_AND2T_59_n95(net373_c1,net373);
INTERCONNECT DFFT_178__FPB_n637_AND2T_55_n91(net374_c1,net374);
INTERCONNECT DFFT_170__FPB_n629_OR2T_47_n83(net375_c1,net375);
INTERCONNECT DFFT_203__FPB_n662_DFFT_204__FPB_n663(net376_c1,net376);
INTERCONNECT DFFT_211__FPB_n670_AND2T_78_n114(net377_c1,net377);
INTERCONNECT DFFT_195__FPB_n654_AND2T_65_n101(net378_c1,net378);
INTERCONNECT DFFT_187__FPB_n646_OR2T_61_n97(net379_c1,net379);
INTERCONNECT DFFT_179__FPB_n638_OR2T_58_n94(net380_c1,net380);
INTERCONNECT DFFT_260__FPB_n719_DFFT_261__FPB_n720(net381_c1,net381);
INTERCONNECT DFFT_204__FPB_n663_DFFT_205__FPB_n664(net382_c1,net382);
INTERCONNECT DFFT_188__FPB_n647_Split_HOLD_869(net383_c1,net383);
INTERCONNECT DFFT_180__FPB_n639_DFFT_181__FPB_n640(net384_c1,net384);
INTERCONNECT DFFT_132__FPB_n591_DFFT_133__FPB_n592(net385_c1,net385);
INTERCONNECT DFFT_212__FPB_n671_OR2T_79_n115(net386_c1,net386);
INTERCONNECT DFFT_196__FPB_n655_Split_HOLD_875(net387_c1,net387);
INTERCONNECT DFFT_205__FPB_n664_DFFT_206__FPB_n665(net388_c1,net388);
INTERCONNECT DFFT_189__FPB_n648_DFFT_190__FPB_n649(net389_c1,net389);
INTERCONNECT DFFT_133__FPB_n592_DFFT_134__FPB_n593(net390_c1,net390);
INTERCONNECT DFFT_221__FPB_n680_AND2T_90_n126(net391_c1,net391);
INTERCONNECT DFFT_213__FPB_n672_OR2T_80_n116(net392_c1,net392);
INTERCONNECT DFFT_197__FPB_n656_OR2T_68_n104(net393_c1,net393);
INTERCONNECT DFFT_222__FPB_n681_Split_HOLD_873(net394_c1,net394);
INTERCONNECT DFFT_190__FPB_n649_DFFT_191__FPB_n650(net395_c1,net395);
INTERCONNECT DFFT_134__FPB_n593_DFFT_135__FPB_n594(net396_c1,net396);
INTERCONNECT DFFT_214__FPB_n673_AND2T_81_n117(net397_c1,net397);
INTERCONNECT DFFT_206__FPB_n665_AND2T_72_n108(net398_c1,net398);
INTERCONNECT DFFT_198__FPB_n657_OR2T_69_n105(net399_c1,net399);
INTERCONNECT DFFT_223__FPB_n682_DFFT_224__FPB_n683(net400_c1,net400);
INTERCONNECT DFFT_135__FPB_n594_DFFT_136__FPB_n595(net401_c1,net401);
INTERCONNECT DFFT_231__FPB_n690_OR2T_99_n135(net402_c1,net402);
INTERCONNECT DFFT_215__FPB_n674_OR2T_87_n123(net403_c1,net403);
INTERCONNECT DFFT_207__FPB_n666_AND2T_73_n109(net404_c1,net404);
INTERCONNECT DFFT_199__FPB_n658_OR2T_70_n106(net405_c1,net405);
INTERCONNECT DFFT_232__FPB_n691_DFFT_233__FPB_n692(net406_c1,net406);
INTERCONNECT DFFT_216__FPB_n675_DFFT_217__FPB_n676(net407_c1,net407);
INTERCONNECT DFFT_200__FPB_n659_Split_HOLD_874(net408_c1,net408);
INTERCONNECT DFFT_136__FPB_n595_DFFT_137__FPB_n596(net409_c1,net409);
INTERCONNECT DFFT_224__FPB_n683_AND2T_91_n127(net410_c1,net410);
INTERCONNECT DFFT_208__FPB_n667_AND2T_74_n110(net411_c1,net411);
INTERCONNECT DFFT_233__FPB_n692_DFFT_234__FPB_n693(net412_c1,net412);
INTERCONNECT DFFT_225__FPB_n684_DFFT_226__FPB_n685(net413_c1,net413);
INTERCONNECT DFFT_217__FPB_n676_DFFT_218__FPB_n677(net414_c1,net414);
INTERCONNECT DFFT_137__FPB_n596_DFFT_121__FBL_n580(net415_c1,net415);
INTERCONNECT DFFT_209__FPB_n668_AND2T_76_n112(net416_c1,net416);
INTERCONNECT DFFT_234__FPB_n693_DFFT_235__FPB_n694(net417_c1,net417);
INTERCONNECT DFFT_218__FPB_n677_DFFT_219__FPB_n678(net418_c1,net418);
INTERCONNECT DFFT_138__FPB_n597_DFFT_139__FPB_n598(net419_c1,net419);
INTERCONNECT DFFT_226__FPB_n685_Split_HOLD_876(net420_c1,net420);
INTERCONNECT DFFT_210__FPB_n669_AND2T_77_n113(net421_c1,net421);
INTERCONNECT DFFT_235__FPB_n694_DFFT_236__FPB_n695(net422_c1,net422);
INTERCONNECT DFFT_227__FPB_n686_DFFT_228__FPB_n687(net423_c1,net423);
INTERCONNECT DFFT_219__FPB_n678_DFFT_220__FPB_n679(net424_c1,net424);
INTERCONNECT DFFT_139__FPB_n598_DFFT_140__FPB_n599(net425_c1,net425);
INTERCONNECT DFFT_236__FPB_n695_Split_HOLD_870(net426_c1,net426);
INTERCONNECT DFFT_220__FPB_n679_DFFT_221__FPB_n680(net427_c1,net427);
INTERCONNECT DFFT_140__FPB_n599_DFFT_122__FBL_n581(net428_c1,net428);
INTERCONNECT DFFT_228__FPB_n687_AND2T_93_n129(net429_c1,net429);
INTERCONNECT DFFT_237__FPB_n696_AND2T_100_n136(net430_c1,net430);
INTERCONNECT DFFT_229__FPB_n688_AND2T_94_n130(net431_c1,net431);
INTERCONNECT DFFT_238__FPB_n697_AND2T_108_n150(net432_c1,net432);
INTERCONNECT DFFT_230__FPB_n689_OR2T_98_n134(net433_c1,net433);
INTERCONNECT DFFT_239__FPB_n698_AND2T_109_n151(net434_c1,net434);
INTERCONNECT DFFT_240__FPB_n699_DFFT_241__FPB_n700(net435_c1,net435);
INTERCONNECT DFFT_245_state_obs0_state_obs0_Pad(net436_c1,state_obs0_Pad);
INTERCONNECT DFFT_251_state_obs1_state_obs1_Pad(net437_c1,state_obs1_Pad);
INTERCONNECT DFFT_259_state_obs2_state_obs2_Pad(net438_c1,state_obs2_Pad);
INTERCONNECT DFFT_267_state_obs3_state_obs3_Pad(net439_c1,state_obs3_Pad);
INTERCONNECT DFFT_105_state0_buf_DFFT_119__PIPL_n170(net440_c1,net440);
INTERCONNECT DFFT_106_state1_buf_DFFT_120__PIPL_n171(net441_c1,net441);
INTERCONNECT SplitCLK_0_771_SplitCLK_0_389(net442_c1,net442);
INTERCONNECT SplitCLK_0_771_SplitCLK_2_518(net443_c1,net443);
INTERCONNECT SplitCLK_4_770_DFFT_198__FPB_n657(net444_c1,net444);
INTERCONNECT SplitCLK_2_769_DFFT_189__FPB_n648(net445_c1,net445);
INTERCONNECT SplitCLK_4_768_DFFT_197__FPB_n656(net446_c1,net446);
INTERCONNECT SplitCLK_2_767_DFFT_188__FPB_n647(net447_c1,net447);
INTERCONNECT SplitCLK_4_766_DFFT_196__FPB_n655(net448_c1,net448);
INTERCONNECT SplitCLK_4_765_DFFT_179__FPB_n638(net449_c1,net449);
INTERCONNECT SplitCLK_2_764_DFFT_187__FPB_n646(net450_c1,net450);
INTERCONNECT SplitCLK_2_763_DFFT_195__FPB_n654(net451_c1,net451);
INTERCONNECT SplitCLK_4_762_DFFT_178__FPB_n637(net452_c1,net452);
INTERCONNECT SplitCLK_4_761_DFFT_186__FPB_n645(net453_c1,net453);
INTERCONNECT SplitCLK_4_760_DFFT_194__FPB_n653(net454_c1,net454);
INTERCONNECT SplitCLK_2_759_DFFT_258__FPB_n717(net455_c1,net455);
INTERCONNECT SplitCLK_4_758_DFFT_266__FPB_n725(net456_c1,net456);
INTERCONNECT SplitCLK_2_757_DFFT_169__FPB_n628(net457_c1,net457);
INTERCONNECT SplitCLK_4_756_DFFT_177__FPB_n636(net458_c1,net458);
INTERCONNECT SplitCLK_2_755_DFFT_185__FPB_n644(net459_c1,net459);
INTERCONNECT SplitCLK_2_754_DFFT_193__FPB_n652(net460_c1,net460);
INTERCONNECT SplitCLK_4_753_DFFT_249__FPB_n708(net461_c1,net461);
INTERCONNECT SplitCLK_2_752_DFFT_265__FPB_n724(net462_c1,net462);
INTERCONNECT SplitCLK_4_751_DFFT_168__FPB_n627(net463_c1,net463);
INTERCONNECT SplitCLK_4_750_DFFT_176__FPB_n635(net464_c1,net464);
INTERCONNECT SplitCLK_4_749_DFFT_184__FPB_n643(net465_c1,net465);
INTERCONNECT SplitCLK_2_748_DFFT_192__FPB_n651(net466_c1,net466);
INTERCONNECT SplitCLK_2_747_DFFT_248__FPB_n707(net467_c1,net467);
INTERCONNECT SplitCLK_2_746_DFFT_264__FPB_n723(net468_c1,net468);
INTERCONNECT SplitCLK_2_745_NOTT_112_n160(net469_c1,net469);
INTERCONNECT SplitCLK_4_744_NOTT_111_n153(net470_c1,net470);
INTERCONNECT SplitCLK_2_743_DFFT_239__FPB_n698(net471_c1,net471);
INTERCONNECT SplitCLK_2_742_DFFT_159__FPB_n618(net472_c1,net472);
INTERCONNECT SplitCLK_4_741_DFFT_167__FPB_n626(net473_c1,net473);
INTERCONNECT SplitCLK_4_740_DFFT_175__FPB_n634(net474_c1,net474);
INTERCONNECT SplitCLK_2_739_DFFT_183__FPB_n642(net475_c1,net475);
INTERCONNECT SplitCLK_2_738_DFFT_191__FPB_n650(net476_c1,net476);
INTERCONNECT SplitCLK_4_737_DFFT_247__FPB_n706(net477_c1,net477);
INTERCONNECT SplitCLK_2_736_DFFT_255__FPB_n714(net478_c1,net478);
INTERCONNECT SplitCLK_4_735_DFFT_238__FPB_n697(net479_c1,net479);
INTERCONNECT SplitCLK_4_734_DFFT_190__FPB_n649(net480_c1,net480);
INTERCONNECT SplitCLK_4_733_DFFT_158__FPB_n617(net481_c1,net481);
INTERCONNECT SplitCLK_2_732_DFFT_174__FPB_n633(net482_c1,net482);
INTERCONNECT SplitCLK_4_731_DFFT_182__FPB_n641(net483_c1,net483);
INTERCONNECT SplitCLK_4_730_DFFT_246__FPB_n705(net484_c1,net484);
INTERCONNECT SplitCLK_4_729_DFFT_254__FPB_n713(net485_c1,net485);
INTERCONNECT SplitCLK_2_728_DFFT_229__FPB_n688(net486_c1,net486);
INTERCONNECT SplitCLK_2_727_DFFT_237__FPB_n696(net487_c1,net487);
INTERCONNECT SplitCLK_4_726_DFFT_149__FPB_n608(net488_c1,net488);
INTERCONNECT SplitCLK_4_725_DFFT_157__FPB_n616(net489_c1,net489);
INTERCONNECT SplitCLK_4_724_DFFT_165__FPB_n624(net490_c1,net490);
INTERCONNECT SplitCLK_4_723_DFFT_173__FPB_n632(net491_c1,net491);
INTERCONNECT SplitCLK_4_722_DFFT_181__FPB_n640(net492_c1,net492);
INTERCONNECT SplitCLK_2_721_DFFT_253__FPB_n712(net493_c1,net493);
INTERCONNECT SplitCLK_4_720_DFFT_261__FPB_n720(net494_c1,net494);
INTERCONNECT SplitCLK_4_719_DFFT_228__FPB_n687(net495_c1,net495);
INTERCONNECT SplitCLK_4_718_DFFT_236__FPB_n695(net496_c1,net496);
INTERCONNECT SplitCLK_4_717_DFFT_180__FPB_n639(net497_c1,net497);
INTERCONNECT SplitCLK_2_716_DFFT_260__FPB_n719(net498_c1,net498);
INTERCONNECT SplitCLK_2_715_DFFT_148__FPB_n607(net499_c1,net499);
INTERCONNECT SplitCLK_2_714_DFFT_156__FPB_n615(net500_c1,net500);
INTERCONNECT SplitCLK_2_713_DFFT_164__FPB_n623(net501_c1,net501);
INTERCONNECT SplitCLK_2_712_DFFT_172__FPB_n631(net502_c1,net502);
INTERCONNECT SplitCLK_2_711_DFFT_244__FPB_n703(net503_c1,net503);
INTERCONNECT SplitCLK_4_710_DFFT_252__FPB_n711(net504_c1,net504);
INTERCONNECT SplitCLK_2_709_DFFT_139__FPB_n598(net505_c1,net505);
INTERCONNECT SplitCLK_4_708_DFFT_219__FPB_n678(net506_c1,net506);
INTERCONNECT SplitCLK_4_707_DFFT_227__FPB_n686(net507_c1,net507);
INTERCONNECT SplitCLK_4_706_DFFT_235__FPB_n694(net508_c1,net508);
INTERCONNECT SplitCLK_4_705_DFFT_147__FPB_n606(net509_c1,net509);
INTERCONNECT SplitCLK_4_704_DFFT_155__FPB_n614(net510_c1,net510);
INTERCONNECT SplitCLK_4_703_DFFT_163__FPB_n622(net511_c1,net511);
INTERCONNECT SplitCLK_2_702_DFFT_171__FPB_n630(net512_c1,net512);
INTERCONNECT SplitCLK_4_701_DFFT_243__FPB_n702(net513_c1,net513);
INTERCONNECT SplitCLK_4_700_DFFT_138__FPB_n597(net514_c1,net514);
INTERCONNECT SplitCLK_4_699_DFFT_218__FPB_n677(net515_c1,net515);
INTERCONNECT SplitCLK_2_698_DFFT_226__FPB_n685(net516_c1,net516);
INTERCONNECT SplitCLK_2_697_DFFT_234__FPB_n693(net517_c1,net517);
INTERCONNECT SplitCLK_2_696_DFFT_170__FPB_n629(net518_c1,net518);
INTERCONNECT SplitCLK_2_695_DFFT_250__FPB_n709(net519_c1,net519);
INTERCONNECT SplitCLK_2_694_DFFT_146__FPB_n605(net520_c1,net520);
INTERCONNECT SplitCLK_4_693_DFFT_154__FPB_n613(net521_c1,net521);
INTERCONNECT SplitCLK_2_692_DFFT_162__FPB_n621(net522_c1,net522);
INTERCONNECT SplitCLK_2_691_DFFT_242__FPB_n701(net523_c1,net523);
INTERCONNECT SplitCLK_2_690_DFFT_137__FPB_n596(net524_c1,net524);
INTERCONNECT SplitCLK_4_689_DFFT_209__FPB_n668(net525_c1,net525);
INTERCONNECT SplitCLK_2_688_DFFT_217__FPB_n676(net526_c1,net526);
INTERCONNECT SplitCLK_2_687_DFFT_225__FPB_n684(net527_c1,net527);
INTERCONNECT SplitCLK_4_686_DFFT_233__FPB_n692(net528_c1,net528);
INTERCONNECT SplitCLK_2_685_DFFT_145__FPB_n604(net529_c1,net529);
INTERCONNECT SplitCLK_2_684_DFFT_153__FPB_n612(net530_c1,net530);
INTERCONNECT SplitCLK_4_683_DFFT_161__FPB_n620(net531_c1,net531);
INTERCONNECT SplitCLK_4_682_DFFT_241__FPB_n700(net532_c1,net532);
INTERCONNECT SplitCLK_2_681_DFFT_129__FBL_n588(net533_c1,net533);
INTERCONNECT SplitCLK_4_680_OR2T_99_n135(net534_c1,net534);
INTERCONNECT SplitCLK_2_679_OR2T_98_n134(net535_c1,net535);
INTERCONNECT SplitCLK_4_678_OR2T_89_n125(net536_c1,net536);
INTERCONNECT SplitCLK_2_677_OR2T_97_n133(net537_c1,net537);
INTERCONNECT SplitCLK_4_676_OR2T_88_n124(net538_c1,net538);
INTERCONNECT SplitCLK_4_675_OR2T_96_n132(net539_c1,net539);
INTERCONNECT SplitCLK_2_674_DFFT_240__FPB_n699(net540_c1,net540);
INTERCONNECT SplitCLK_4_673_OR2T_79_n115(net541_c1,net541);
INTERCONNECT SplitCLK_2_672_OR2T_87_n123(net542_c1,net542);
INTERCONNECT SplitCLK_2_671_OR2T_95_n131(net543_c1,net543);
INTERCONNECT SplitCLK_4_670_DFFT_136__FPB_n595(net544_c1,net544);
INTERCONNECT SplitCLK_2_669_DFFT_208__FPB_n667(net545_c1,net545);
INTERCONNECT SplitCLK_4_668_DFFT_216__FPB_n675(net546_c1,net546);
INTERCONNECT SplitCLK_2_667_DFFT_224__FPB_n683(net547_c1,net547);
INTERCONNECT SplitCLK_2_666_DFFT_232__FPB_n691(net548_c1,net548);
INTERCONNECT SplitCLK_2_665_DFFT_160__FPB_n619(net549_c1,net549);
INTERCONNECT SplitCLK_4_664_DFFT_144__FPB_n603(net550_c1,net550);
INTERCONNECT SplitCLK_2_663_DFFT_152__FPB_n611(net551_c1,net551);
INTERCONNECT SplitCLK_4_662_OR2T_69_n105(net552_c1,net552);
INTERCONNECT SplitCLK_2_661_OR2T_68_n104(net553_c1,net553);
INTERCONNECT SplitCLK_4_660_OR2T_84_n120(net554_c1,net554);
INTERCONNECT SplitCLK_2_659_OR2T_83_n119(net555_c1,net555);
INTERCONNECT SplitCLK_2_658_OR2T_80_n116(net556_c1,net556);
INTERCONNECT SplitCLK_2_657_OR2T_64_n100(net557_c1,net557);
INTERCONNECT SplitCLK_2_656_OR2T_71_n107(net558_c1,net558);
INTERCONNECT SplitCLK_4_655_OR2T_70_n106(net559_c1,net559);
INTERCONNECT SplitCLK_2_654_DFFT_128__FBL_n587(net560_c1,net560);
INTERCONNECT SplitCLK_4_653_DFFT_135__FPB_n594(net561_c1,net561);
INTERCONNECT SplitCLK_2_652_DFFT_207__FPB_n666(net562_c1,net562);
INTERCONNECT SplitCLK_4_651_DFFT_215__FPB_n674(net563_c1,net563);
INTERCONNECT SplitCLK_2_650_DFFT_223__FPB_n682(net564_c1,net564);
INTERCONNECT SplitCLK_4_649_DFFT_231__FPB_n690(net565_c1,net565);
INTERCONNECT SplitCLK_2_648_DFFT_143__FPB_n602(net566_c1,net566);
INTERCONNECT SplitCLK_4_647_DFFT_151__FPB_n610(net567_c1,net567);
INTERCONNECT SplitCLK_2_646_DFFT_127__FBL_n586(net568_c1,net568);
INTERCONNECT SplitCLK_4_645_DFFT_230__FPB_n689(net569_c1,net569);
INTERCONNECT SplitCLK_4_644_DFFT_134__FPB_n593(net570_c1,net570);
INTERCONNECT SplitCLK_4_643_DFFT_206__FPB_n665(net571_c1,net571);
INTERCONNECT SplitCLK_2_642_DFFT_214__FPB_n673(net572_c1,net572);
INTERCONNECT SplitCLK_4_641_DFFT_222__FPB_n681(net573_c1,net573);
INTERCONNECT SplitCLK_2_640_DFFT_150__FPB_n609(net574_c1,net574);
INTERCONNECT SplitCLK_4_639_DFFT_142__FPB_n601(net575_c1,net575);
INTERCONNECT SplitCLK_2_638_DFFT_126__FBL_n585(net576_c1,net576);
INTERCONNECT SplitCLK_2_637_DFFT_133__FPB_n592(net577_c1,net577);
INTERCONNECT SplitCLK_4_636_DFFT_205__FPB_n664(net578_c1,net578);
INTERCONNECT SplitCLK_2_635_DFFT_213__FPB_n672(net579_c1,net579);
INTERCONNECT SplitCLK_4_634_DFFT_221__FPB_n680(net580_c1,net580);
INTERCONNECT SplitCLK_4_633_DFFT_141__FPB_n600(net581_c1,net581);
INTERCONNECT SplitCLK_2_632_DFFT_125__FBL_n584(net582_c1,net582);
INTERCONNECT SplitCLK_4_631_DFFT_140__FPB_n599(net583_c1,net583);
INTERCONNECT SplitCLK_4_630_DFFT_220__FPB_n679(net584_c1,net584);
INTERCONNECT SplitCLK_4_629_DFFT_132__FPB_n591(net585_c1,net585);
INTERCONNECT SplitCLK_2_628_DFFT_204__FPB_n663(net586_c1,net586);
INTERCONNECT SplitCLK_2_627_DFFT_212__FPB_n671(net587_c1,net587);
INTERCONNECT SplitCLK_4_626_DFFT_124__FBL_n583(net588_c1,net588);
INTERCONNECT SplitCLK_4_625_DFFT_203__FPB_n662(net589_c1,net589);
INTERCONNECT SplitCLK_2_624_DFFT_211__FPB_n670(net590_c1,net590);
INTERCONNECT SplitCLK_4_623_DFFT_123__FBL_n582(net591_c1,net591);
INTERCONNECT SplitCLK_2_622_DFFT_131__FBL_n590(net592_c1,net592);
INTERCONNECT SplitCLK_2_621_DFFT_210__FPB_n669(net593_c1,net593);
INTERCONNECT SplitCLK_4_620_DFFT_202__FPB_n661(net594_c1,net594);
INTERCONNECT SplitCLK_2_619_DFFT_114__FPB_n165(net595_c1,net595);
INTERCONNECT SplitCLK_4_618_DFFT_130__FBL_n589(net596_c1,net596);
INTERCONNECT SplitCLK_4_617_DFFT_122__FBL_n581(net597_c1,net597);
INTERCONNECT SplitCLK_4_616_DFFT_201__FPB_n660(net598_c1,net598);
INTERCONNECT SplitCLK_4_615_DFFT_113__FPB_n164(net599_c1,net599);
INTERCONNECT SplitCLK_4_614_DFFT_121__FBL_n580(net600_c1,net600);
INTERCONNECT SplitCLK_2_613_DFFT_200__FPB_n659(net601_c1,net601);
INTERCONNECT SplitCLK_2_612_AND2T_78_n114(net602_c1,net602);
INTERCONNECT SplitCLK_2_611_AND2T_86_n122(net603_c1,net603);
INTERCONNECT SplitCLK_4_610_AND2T_94_n130(net604_c1,net604);
INTERCONNECT SplitCLK_2_609_AND2T_93_n129(net605_c1,net605);
INTERCONNECT SplitCLK_2_608_AND2T_85_n121(net606_c1,net606);
INTERCONNECT SplitCLK_4_607_AND2T_92_n128(net607_c1,net607);
INTERCONNECT SplitCLK_2_606_AND2T_91_n127(net608_c1,net608);
INTERCONNECT SplitCLK_2_605_AND2T_67_n103(net609_c1,net609);
INTERCONNECT SplitCLK_4_604_AND2T_82_n118(net610_c1,net610);
INTERCONNECT SplitCLK_4_603_AND2T_90_n126(net611_c1,net611);
INTERCONNECT SplitCLK_4_602_AND2T_66_n102(net612_c1,net612);
INTERCONNECT SplitCLK_4_601_AND2T_74_n110(net613_c1,net613);
INTERCONNECT SplitCLK_4_600_AND2T_73_n109(net614_c1,net614);
INTERCONNECT SplitCLK_2_599_AND2T_81_n117(net615_c1,net615);
INTERCONNECT SplitCLK_4_598_AND2T_65_n101(net616_c1,net616);
INTERCONNECT SplitCLK_4_597_AND2T_72_n108(net617_c1,net617);
INTERCONNECT SplitCLK_2_596_DFFT_119__PIPL_n170(net618_c1,net618);
INTERCONNECT SplitCLK_4_595_DFFT_118__PIPL_n169(net619_c1,net619);
INTERCONNECT SplitCLK_4_594_DFFT_117__PIPL_n168(net620_c1,net620);
INTERCONNECT SplitCLK_4_593_NOTT_26_n62(net621_c1,net621);
INTERCONNECT SplitCLK_2_592_NOTT_25_n61(net622_c1,net622);
INTERCONNECT SplitCLK_2_591_NOTT_16_n52(net623_c1,net623);
INTERCONNECT SplitCLK_4_590_NOTT_24_n60(net624_c1,net624);
INTERCONNECT SplitCLK_4_589_NOTT_23_n59(net625_c1,net625);
INTERCONNECT SplitCLK_4_588_NOTT_14_n50(net626_c1,net626);
INTERCONNECT SplitCLK_4_587_NOTT_12_n48(net627_c1,net627);
INTERCONNECT SplitCLK_4_586_NOTT_10_n46(net628_c1,net628);
INTERCONNECT SplitCLK_2_585_DFFT_116__PIPL_n167(net629_c1,net629);
INTERCONNECT SplitCLK_4_584_DFFT_115__PIPL_n166(net630_c1,net630);
INTERCONNECT SplitCLK_4_583_OR2T_58_n94(net631_c1,net631);
INTERCONNECT SplitCLK_2_582_OR2T_57_n93(net632_c1,net632);
INTERCONNECT SplitCLK_2_581_OR2T_56_n92(net633_c1,net633);
INTERCONNECT SplitCLK_2_580_OR2T_47_n83(net634_c1,net634);
INTERCONNECT SplitCLK_4_579_OR2T_46_n82(net635_c1,net635);
INTERCONNECT SplitCLK_4_578_OR2T_54_n90(net636_c1,net636);
INTERCONNECT SplitCLK_2_577_OR2T_61_n97(net637_c1,net637);
INTERCONNECT SplitCLK_4_576_OR2T_45_n81(net638_c1,net638);
INTERCONNECT SplitCLK_2_575_OR2T_60_n96(net639_c1,net639);
INTERCONNECT SplitCLK_4_574_OR2T_50_n86(net640_c1,net640);
INTERCONNECT SplitCLK_4_573_OR2T_34_n70(net641_c1,net641);
INTERCONNECT SplitCLK_2_572_OR2T_33_n69(net642_c1,net642);
INTERCONNECT SplitCLK_2_571_OR2T_40_n76(net643_c1,net643);
INTERCONNECT SplitCLK_2_570_OR2T_22_n58(net644_c1,net644);
INTERCONNECT SplitCLK_2_569_OR2T_21_n57(net645_c1,net645);
INTERCONNECT SplitCLK_2_568_OR2T_11_n47(net646_c1,net646);
INTERCONNECT SplitCLK_2_567_DFFT_120__PIPL_n171(net647_c1,net647);
INTERCONNECT SplitCLK_2_566_DFFT_267_state_obs3(net648_c1,net648);
INTERCONNECT SplitCLK_2_565_DFFT_259_state_obs2(net649_c1,net649);
INTERCONNECT SplitCLK_4_564_AND2T_59_n95(net650_c1,net650);
INTERCONNECT SplitCLK_2_563_AND2T_49_n85(net651_c1,net651);
INTERCONNECT SplitCLK_2_562_AND2T_48_n84(net652_c1,net652);
INTERCONNECT SplitCLK_4_561_AND2T_63_n99(net653_c1,net653);
INTERCONNECT SplitCLK_2_560_AND2T_39_n75(net654_c1,net654);
INTERCONNECT SplitCLK_4_559_AND2T_55_n91(net655_c1,net655);
INTERCONNECT SplitCLK_4_558_AND2T_62_n98(net656_c1,net656);
INTERCONNECT SplitCLK_4_557_AND2T_53_n89(net657_c1,net657);
INTERCONNECT SplitCLK_2_556_AND2T_29_n65(net658_c1,net658);
INTERCONNECT SplitCLK_4_555_AND2T_37_n73(net659_c1,net659);
INTERCONNECT SplitCLK_4_554_AND2T_52_n88(net660_c1,net660);
INTERCONNECT SplitCLK_2_553_AND2T_28_n64(net661_c1,net661);
INTERCONNECT SplitCLK_4_552_AND2T_36_n72(net662_c1,net662);
INTERCONNECT SplitCLK_2_551_AND2T_44_n80(net663_c1,net663);
INTERCONNECT SplitCLK_2_550_AND2T_43_n79(net664_c1,net664);
INTERCONNECT SplitCLK_2_549_AND2T_51_n87(net665_c1,net665);
INTERCONNECT SplitCLK_2_548_AND2T_19_n55(net666_c1,net666);
INTERCONNECT SplitCLK_4_547_AND2T_27_n63(net667_c1,net667);
INTERCONNECT SplitCLK_4_546_AND2T_35_n71(net668_c1,net668);
INTERCONNECT SplitCLK_2_545_AND2T_42_n78(net669_c1,net669);
INTERCONNECT SplitCLK_4_544_AND2T_18_n54(net670_c1,net670);
INTERCONNECT SplitCLK_4_543_AND2T_41_n77(net671_c1,net671);
INTERCONNECT SplitCLK_2_542_AND2T_17_n53(net672_c1,net672);
INTERCONNECT SplitCLK_4_541_AND2T_32_n68(net673_c1,net673);
INTERCONNECT SplitCLK_2_540_AND2T_31_n67(net674_c1,net674);
INTERCONNECT SplitCLK_4_539_AND2T_15_n51(net675_c1,net675);
INTERCONNECT SplitCLK_2_538_AND2T_30_n66(net676_c1,net676);
INTERCONNECT SplitCLK_2_537_AND2T_13_n49(net677_c1,net677);
INTERCONNECT SplitCLK_2_536_AND2T_20_n56(net678_c1,net678);
INTERCONNECT SplitCLK_2_535_XOR2T_75_n111(net679_c1,net679);
INTERCONNECT SplitCLK_4_534_NOTT_9_n45(net680_c1,net680);
INTERCONNECT SplitCLK_4_533_DFFT_106_state1_buf(net681_c1,net681);
INTERCONNECT SplitCLK_4_532_AND2T_8_n44(net682_c1,net682);
INTERCONNECT SplitCLK_2_531_DFFT_104_state_obs3_buf(net683_c1,net683);
INTERCONNECT SplitCLK_2_530_DFFT_103_state_obs2_buf(net684_c1,net684);
INTERCONNECT SplitCLK_4_529_DFFT_102_state_obs1_buf(net685_c1,net685);
INTERCONNECT SplitCLK_2_528_DFFT_101_state_obs0_buf(net686_c1,net686);
INTERCONNECT SplitCLK_4_527_AND2T_109_n151(net687_c1,net687);
INTERCONNECT SplitCLK_2_526_AND2T_108_n150(net688_c1,net688);
INTERCONNECT SplitCLK_2_525_AND2T_107_n149(net689_c1,net689);
INTERCONNECT SplitCLK_2_524_AND2T_110_n152(net690_c1,net690);
INTERCONNECT SplitCLK_4_523_AND2T_100_n136(net691_c1,net691);
INTERCONNECT SplitCLK_2_522_DFFT_245_state_obs0(net692_c1,net692);
INTERCONNECT SplitCLK_2_521_DFFT_251_state_obs1(net693_c1,net693);
INTERCONNECT SplitCLK_4_520_DFFT_105_state0_buf(net694_c1,net694);
INTERCONNECT SplitCLK_2_519_DFFT_199__FPB_n658(net695_c1,net695);
INTERCONNECT SplitCLK_2_518_SplitCLK_6_453(net696_c1,net696);
INTERCONNECT SplitCLK_2_518_SplitCLK_4_517(net697_c1,net697);
INTERCONNECT SplitCLK_4_517_SplitCLK_0_485(net698_c1,net698);
INTERCONNECT SplitCLK_4_517_SplitCLK_4_516(net699_c1,net699);
INTERCONNECT SplitCLK_4_516_SplitCLK_6_500(net700_c1,net700);
INTERCONNECT SplitCLK_4_516_SplitCLK_4_515(net701_c1,net701);
INTERCONNECT SplitCLK_4_515_SplitCLK_4_507(net702_c1,net702);
INTERCONNECT SplitCLK_4_515_SplitCLK_2_514(net703_c1,net703);
INTERCONNECT SplitCLK_2_514_SplitCLK_6_510(net704_c1,net704);
INTERCONNECT SplitCLK_2_514_SplitCLK_4_513(net705_c1,net705);
INTERCONNECT SplitCLK_4_513_SplitCLK_4_511(net706_c1,net706);
INTERCONNECT SplitCLK_4_513_SplitCLK_6_512(net707_c1,net707);
INTERCONNECT SplitCLK_6_512_SplitCLK_4_749(net708_c1,net708);
INTERCONNECT SplitCLK_6_512_SplitCLK_2_755(net709_c1,net709);
INTERCONNECT SplitCLK_4_511_SplitCLK_4_731(net710_c1,net710);
INTERCONNECT SplitCLK_4_511_SplitCLK_2_739(net711_c1,net711);
INTERCONNECT SplitCLK_6_510_SplitCLK_0_508(net712_c1,net712);
INTERCONNECT SplitCLK_6_510_SplitCLK_2_509(net713_c1,net713);
INTERCONNECT SplitCLK_2_509_SplitCLK_2_687(net714_c1,net714);
INTERCONNECT SplitCLK_2_509_SplitCLK_4_761(net715_c1,net715);
INTERCONNECT SplitCLK_0_508_SplitCLK_4_641(net716_c1,net716);
INTERCONNECT SplitCLK_0_508_SplitCLK_2_698(net717_c1,net717);
INTERCONNECT SplitCLK_4_507_SplitCLK_4_503(net718_c1,net718);
INTERCONNECT SplitCLK_4_507_SplitCLK_4_506(net719_c1,net719);
INTERCONNECT SplitCLK_4_506_SplitCLK_4_504(net720_c1,net720);
INTERCONNECT SplitCLK_4_506_SplitCLK_2_505(net721_c1,net721);
INTERCONNECT SplitCLK_2_505_SplitCLK_2_619(net722_c1,net722);
INTERCONNECT SplitCLK_2_505_SplitCLK_4_722(net723_c1,net723);
INTERCONNECT SplitCLK_4_504_SplitCLK_4_625(net724_c1,net724);
INTERCONNECT SplitCLK_4_504_SplitCLK_2_628(net725_c1,net725);
INTERCONNECT SplitCLK_4_503_SplitCLK_0_501(net726_c1,net726);
INTERCONNECT SplitCLK_4_503_SplitCLK_6_502(net727_c1,net727);
INTERCONNECT SplitCLK_6_502_SplitCLK_4_636(net728_c1,net728);
INTERCONNECT SplitCLK_6_502_SplitCLK_2_650(net729_c1,net729);
INTERCONNECT SplitCLK_0_501_SplitCLK_4_643(net730_c1,net730);
INTERCONNECT SplitCLK_0_501_SplitCLK_2_667(net731_c1,net731);
INTERCONNECT SplitCLK_6_500_SplitCLK_0_492(net732_c1,net732);
INTERCONNECT SplitCLK_6_500_SplitCLK_2_499(net733_c1,net733);
INTERCONNECT SplitCLK_2_499_SplitCLK_2_495(net734_c1,net734);
INTERCONNECT SplitCLK_2_499_SplitCLK_4_498(net735_c1,net735);
INTERCONNECT SplitCLK_4_498_SplitCLK_0_496(net736_c1,net736);
INTERCONNECT SplitCLK_4_498_SplitCLK_6_497(net737_c1,net737);
INTERCONNECT SplitCLK_6_497_SplitCLK_4_564(net738_c1,net738);
INTERCONNECT SplitCLK_6_497_SplitCLK_2_624(net739_c1,net739);
INTERCONNECT SplitCLK_0_496_SplitCLK_2_612(net740_c1,net740);
INTERCONNECT SplitCLK_0_496_SplitCLK_4_623(net741_c1,net741);
INTERCONNECT SplitCLK_2_495_SplitCLK_0_493(net742_c1,net742);
INTERCONNECT SplitCLK_2_495_SplitCLK_4_494(net743_c1,net743);
INTERCONNECT SplitCLK_4_494_SplitCLK_2_608(net744_c1,net744);
INTERCONNECT SplitCLK_4_494_SplitCLK_2_646(net745_c1,net745);
INTERCONNECT SplitCLK_0_493_SplitCLK_2_592(net746_c1,net746);
INTERCONNECT SplitCLK_0_493_SplitCLK_4_626(net747_c1,net747);
INTERCONNECT SplitCLK_0_492_SplitCLK_6_488(net748_c1,net748);
INTERCONNECT SplitCLK_0_492_SplitCLK_4_491(net749_c1,net749);
INTERCONNECT SplitCLK_4_491_SplitCLK_0_489(net750_c1,net750);
INTERCONNECT SplitCLK_4_491_SplitCLK_2_490(net751_c1,net751);
INTERCONNECT SplitCLK_2_490_SplitCLK_4_607(net752_c1,net752);
INTERCONNECT SplitCLK_2_490_SplitCLK_2_677(net753_c1,net753);
INTERCONNECT SplitCLK_0_489_SplitCLK_4_645(net754_c1,net754);
INTERCONNECT SplitCLK_0_489_SplitCLK_4_770(net755_c1,net755);
INTERCONNECT SplitCLK_6_488_SplitCLK_0_486(net756_c1,net756);
INTERCONNECT SplitCLK_6_488_SplitCLK_6_487(net757_c1,net757);
INTERCONNECT SplitCLK_6_487_SplitCLK_2_556(net758_c1,net758);
INTERCONNECT SplitCLK_6_487_SplitCLK_4_719(net759_c1,net759);
INTERCONNECT SplitCLK_0_486_SplitCLK_4_675(net760_c1,net760);
INTERCONNECT SplitCLK_0_486_SplitCLK_4_707(net761_c1,net761);
INTERCONNECT SplitCLK_0_485_SplitCLK_6_469(net762_c1,net762);
INTERCONNECT SplitCLK_0_485_SplitCLK_4_484(net763_c1,net763);
INTERCONNECT SplitCLK_4_484_SplitCLK_4_476(net764_c1,net764);
INTERCONNECT SplitCLK_4_484_SplitCLK_2_483(net765_c1,net765);
INTERCONNECT SplitCLK_2_483_SplitCLK_6_479(net766_c1,net766);
INTERCONNECT SplitCLK_2_483_SplitCLK_4_482(net767_c1,net767);
INTERCONNECT SplitCLK_4_482_SplitCLK_0_480(net768_c1,net768);
INTERCONNECT SplitCLK_4_482_SplitCLK_6_481(net769_c1,net769);
INTERCONNECT SplitCLK_6_481_SplitCLK_4_620(net770_c1,net770);
INTERCONNECT SplitCLK_6_481_SplitCLK_4_744(net771_c1,net771);
INTERCONNECT SplitCLK_0_480_SplitCLK_4_615(net772_c1,net772);
INTERCONNECT SplitCLK_0_480_SplitCLK_4_616(net773_c1,net773);
INTERCONNECT SplitCLK_6_479_SplitCLK_0_477(net774_c1,net774);
INTERCONNECT SplitCLK_6_479_SplitCLK_2_478(net775_c1,net775);
INTERCONNECT SplitCLK_2_478_SplitCLK_4_597(net776_c1,net776);
INTERCONNECT SplitCLK_2_478_SplitCLK_2_679(net777_c1,net777);
INTERCONNECT SplitCLK_0_477_SplitCLK_4_523(net778_c1,net778);
INTERCONNECT SplitCLK_0_477_SplitCLK_4_649(net779_c1,net779);
INTERCONNECT SplitCLK_4_476_SplitCLK_6_472(net780_c1,net780);
INTERCONNECT SplitCLK_4_476_SplitCLK_4_475(net781_c1,net781);
INTERCONNECT SplitCLK_4_475_SplitCLK_0_473(net782_c1,net782);
INTERCONNECT SplitCLK_4_475_SplitCLK_6_474(net783_c1,net783);
INTERCONNECT SplitCLK_6_474_SplitCLK_2_613(net784_c1,net784);
INTERCONNECT SplitCLK_6_474_SplitCLK_4_717(net785_c1,net785);
INTERCONNECT SplitCLK_0_473_SplitCLK_4_630(net786_c1,net786);
INTERCONNECT SplitCLK_0_473_SplitCLK_2_712(net787_c1,net787);
INTERCONNECT SplitCLK_6_472_SplitCLK_4_470(net788_c1,net788);
INTERCONNECT SplitCLK_6_472_SplitCLK_6_471(net789_c1,net789);
INTERCONNECT SplitCLK_6_471_SplitCLK_2_606(net790_c1,net790);
INTERCONNECT SplitCLK_6_471_SplitCLK_4_723(net791_c1,net791);
INTERCONNECT SplitCLK_4_470_SplitCLK_4_558(net792_c1,net792);
INTERCONNECT SplitCLK_4_470_SplitCLK_2_732(net793_c1,net793);
INTERCONNECT SplitCLK_6_469_SplitCLK_4_461(net794_c1,net794);
INTERCONNECT SplitCLK_6_469_SplitCLK_2_468(net795_c1,net795);
INTERCONNECT SplitCLK_2_468_SplitCLK_2_464(net796_c1,net796);
INTERCONNECT SplitCLK_2_468_SplitCLK_4_467(net797_c1,net797);
INTERCONNECT SplitCLK_4_467_SplitCLK_4_465(net798_c1,net798);
INTERCONNECT SplitCLK_4_467_SplitCLK_2_466(net799_c1,net799);
INTERCONNECT SplitCLK_2_466_SplitCLK_2_642(net800_c1,net800);
INTERCONNECT SplitCLK_2_466_SplitCLK_4_680(net801_c1,net801);
INTERCONNECT SplitCLK_4_465_SplitCLK_2_599(net802_c1,net802);
INTERCONNECT SplitCLK_4_465_SplitCLK_2_659(net803_c1,net803);
INTERCONNECT SplitCLK_2_464_SplitCLK_0_462(net804_c1,net804);
INTERCONNECT SplitCLK_2_464_SplitCLK_4_463(net805_c1,net805);
INTERCONNECT SplitCLK_4_463_SplitCLK_2_609(net806_c1,net806);
INTERCONNECT SplitCLK_4_463_SplitCLK_2_671(net807_c1,net807);
INTERCONNECT SplitCLK_0_462_SplitCLK_4_604(net808_c1,net808);
INTERCONNECT SplitCLK_0_462_SplitCLK_2_611(net809_c1,net809);
INTERCONNECT SplitCLK_4_461_SplitCLK_2_457(net810_c1,net810);
INTERCONNECT SplitCLK_4_461_SplitCLK_4_460(net811_c1,net811);
INTERCONNECT SplitCLK_4_460_SplitCLK_0_458(net812_c1,net812);
INTERCONNECT SplitCLK_4_460_SplitCLK_2_459(net813_c1,net813);
INTERCONNECT SplitCLK_2_459_SplitCLK_2_545(net814_c1,net814);
INTERCONNECT SplitCLK_2_459_SplitCLK_4_590(net815_c1,net815);
INTERCONNECT SplitCLK_0_458_SplitCLK_2_605(net816_c1,net816);
INTERCONNECT SplitCLK_0_458_SplitCLK_4_751(net817_c1,net817);
INTERCONNECT SplitCLK_2_457_SplitCLK_0_455(net818_c1,net818);
INTERCONNECT SplitCLK_2_457_SplitCLK_6_456(net819_c1,net819);
INTERCONNECT SplitCLK_6_456_SplitCLK_2_627(net820_c1,net820);
INTERCONNECT SplitCLK_6_456_SplitCLK_4_673(net821_c1,net821);
INTERCONNECT SplitCLK_0_455_SplitCLK_4_766(net822_c1,net822);
INTERCONNECT SplitCLK_0_455_SplitCLK_0_454(net823_c1,net823);
INTERCONNECT SplitCLK_0_454_AND2T_76_n112(net824_c1,net824);
INTERCONNECT SplitCLK_0_454_AND2T_77_n113(net825_c1,net825);
INTERCONNECT SplitCLK_6_453_SplitCLK_0_421(net826_c1,net826);
INTERCONNECT SplitCLK_6_453_SplitCLK_2_452(net827_c1,net827);
INTERCONNECT SplitCLK_2_452_SplitCLK_6_436(net828_c1,net828);
INTERCONNECT SplitCLK_2_452_SplitCLK_4_451(net829_c1,net829);
INTERCONNECT SplitCLK_4_451_SplitCLK_4_443(net830_c1,net830);
INTERCONNECT SplitCLK_4_451_SplitCLK_2_450(net831_c1,net831);
INTERCONNECT SplitCLK_2_450_SplitCLK_6_446(net832_c1,net832);
INTERCONNECT SplitCLK_2_450_SplitCLK_4_449(net833_c1,net833);
INTERCONNECT SplitCLK_4_449_SplitCLK_4_447(net834_c1,net834);
INTERCONNECT SplitCLK_4_449_SplitCLK_0_448(net835_c1,net835);
INTERCONNECT SplitCLK_0_448_SplitCLK_2_685(net836_c1,net836);
INTERCONNECT SplitCLK_0_448_SplitCLK_4_725(net837_c1,net837);
INTERCONNECT SplitCLK_4_447_SplitCLK_4_573(net838_c1,net838);
INTERCONNECT SplitCLK_4_447_SplitCLK_2_742(net839_c1,net839);
INTERCONNECT SplitCLK_6_446_SplitCLK_4_444(net840_c1,net840);
INTERCONNECT SplitCLK_6_446_SplitCLK_2_445(net841_c1,net841);
INTERCONNECT SplitCLK_2_445_SplitCLK_4_618(net842_c1,net842);
INTERCONNECT SplitCLK_2_445_SplitCLK_2_745(net843_c1,net843);
INTERCONNECT SplitCLK_4_444_SplitCLK_4_664(net844_c1,net844);
INTERCONNECT SplitCLK_4_444_SplitCLK_2_681(net845_c1,net845);
INTERCONNECT SplitCLK_4_443_SplitCLK_2_439(net846_c1,net846);
INTERCONNECT SplitCLK_4_443_SplitCLK_2_442(net847_c1,net847);
INTERCONNECT SplitCLK_2_442_SplitCLK_4_440(net848_c1,net848);
INTERCONNECT SplitCLK_2_442_SplitCLK_6_441(net849_c1,net849);
INTERCONNECT SplitCLK_6_441_SplitCLK_2_572(net850_c1,net850);
INTERCONNECT SplitCLK_6_441_SplitCLK_2_669(net851_c1,net851);
INTERCONNECT SplitCLK_4_440_SplitCLK_4_593(net852_c1,net852);
INTERCONNECT SplitCLK_4_440_SplitCLK_2_728(net853_c1,net853);
INTERCONNECT SplitCLK_2_439_SplitCLK_0_437(net854_c1,net854);
INTERCONNECT SplitCLK_2_439_SplitCLK_2_438(net855_c1,net855);
INTERCONNECT SplitCLK_2_438_SplitCLK_2_684(net856_c1,net856);
INTERCONNECT SplitCLK_2_438_SplitCLK_2_694(net857_c1,net857);
INTERCONNECT SplitCLK_0_437_SplitCLK_2_622(net858_c1,net858);
INTERCONNECT SplitCLK_0_437_SplitCLK_4_733(net859_c1,net859);
INTERCONNECT SplitCLK_6_436_SplitCLK_4_428(net860_c1,net860);
INTERCONNECT SplitCLK_6_436_SplitCLK_2_435(net861_c1,net861);
INTERCONNECT SplitCLK_2_435_SplitCLK_6_431(net862_c1,net862);
INTERCONNECT SplitCLK_2_435_SplitCLK_4_434(net863_c1,net863);
INTERCONNECT SplitCLK_4_434_SplitCLK_4_432(net864_c1,net864);
INTERCONNECT SplitCLK_4_434_SplitCLK_6_433(net865_c1,net865);
INTERCONNECT SplitCLK_6_433_SplitCLK_4_614(net866_c1,net866);
INTERCONNECT SplitCLK_6_433_SplitCLK_2_674(net867_c1,net867);
INTERCONNECT SplitCLK_4_432_SplitCLK_4_670(net868_c1,net868);
INTERCONNECT SplitCLK_4_432_SplitCLK_2_690(net869_c1,net869);
INTERCONNECT SplitCLK_6_431_SplitCLK_0_429(net870_c1,net870);
INTERCONNECT SplitCLK_6_431_SplitCLK_6_430(net871_c1,net871);
INTERCONNECT SplitCLK_6_430_SplitCLK_2_522(net872_c1,net872);
INTERCONNECT SplitCLK_6_430_SplitCLK_4_682(net873_c1,net873);
INTERCONNECT SplitCLK_0_429_SplitCLK_4_584(net874_c1,net874);
INTERCONNECT SplitCLK_0_429_SplitCLK_2_711(net875_c1,net875);
INTERCONNECT SplitCLK_4_428_SplitCLK_0_424(net876_c1,net876);
INTERCONNECT SplitCLK_4_428_SplitCLK_4_427(net877_c1,net877);
INTERCONNECT SplitCLK_4_427_SplitCLK_0_425(net878_c1,net878);
INTERCONNECT SplitCLK_4_427_SplitCLK_6_426(net879_c1,net879);
INTERCONNECT SplitCLK_6_426_SplitCLK_2_528(net880_c1,net880);
INTERCONNECT SplitCLK_6_426_SplitCLK_4_653(net881_c1,net881);
INTERCONNECT SplitCLK_0_425_SplitCLK_2_596(net882_c1,net882);
INTERCONNECT SplitCLK_0_425_SplitCLK_4_644(net883_c1,net883);
INTERCONNECT SplitCLK_0_424_SplitCLK_0_422(net884_c1,net884);
INTERCONNECT SplitCLK_0_424_SplitCLK_6_423(net885_c1,net885);
INTERCONNECT SplitCLK_6_423_SplitCLK_2_691(net886_c1,net886);
INTERCONNECT SplitCLK_6_423_SplitCLK_4_701(net887_c1,net887);
INTERCONNECT SplitCLK_0_422_SplitCLK_4_520(net888_c1,net888);
INTERCONNECT SplitCLK_0_422_SplitCLK_2_521(net889_c1,net889);
INTERCONNECT SplitCLK_0_421_SplitCLK_6_405(net890_c1,net890);
INTERCONNECT SplitCLK_0_421_SplitCLK_4_420(net891_c1,net891);
INTERCONNECT SplitCLK_4_420_SplitCLK_0_412(net892_c1,net892);
INTERCONNECT SplitCLK_4_420_SplitCLK_4_419(net893_c1,net893);
INTERCONNECT SplitCLK_4_419_SplitCLK_0_415(net894_c1,net894);
INTERCONNECT SplitCLK_4_419_SplitCLK_2_418(net895_c1,net895);
INTERCONNECT SplitCLK_2_418_SplitCLK_0_416(net896_c1,net896);
INTERCONNECT SplitCLK_2_418_SplitCLK_6_417(net897_c1,net897);
INTERCONNECT SplitCLK_6_417_SplitCLK_2_548(net898_c1,net898);
INTERCONNECT SplitCLK_6_417_SplitCLK_4_601(net899_c1,net899);
INTERCONNECT SplitCLK_0_416_SplitCLK_4_610(net900_c1,net900);
INTERCONNECT SplitCLK_0_416_SplitCLK_4_740(net901_c1,net901);
INTERCONNECT SplitCLK_0_415_SplitCLK_0_413(net902_c1,net902);
INTERCONNECT SplitCLK_0_415_SplitCLK_2_414(net903_c1,net903);
INTERCONNECT SplitCLK_2_414_SplitCLK_2_536(net904_c1,net904);
INTERCONNECT SplitCLK_2_414_SplitCLK_4_541(net905_c1,net905);
INTERCONNECT SplitCLK_0_413_SplitCLK_2_535(net906_c1,net906);
INTERCONNECT SplitCLK_0_413_SplitCLK_4_689(net907_c1,net907);
INTERCONNECT SplitCLK_0_412_SplitCLK_6_408(net908_c1,net908);
INTERCONNECT SplitCLK_0_412_SplitCLK_4_411(net909_c1,net909);
INTERCONNECT SplitCLK_4_411_SplitCLK_0_409(net910_c1,net910);
INTERCONNECT SplitCLK_4_411_SplitCLK_4_410(net911_c1,net911);
INTERCONNECT SplitCLK_4_410_SplitCLK_2_538(net912_c1,net912);
INTERCONNECT SplitCLK_4_410_SplitCLK_2_540(net913_c1,net913);
INTERCONNECT SplitCLK_0_409_SplitCLK_4_554(net914_c1,net914);
INTERCONNECT SplitCLK_0_409_SplitCLK_2_632(net915_c1,net915);
INTERCONNECT SplitCLK_6_408_SplitCLK_0_406(net916_c1,net916);
INTERCONNECT SplitCLK_6_408_SplitCLK_2_407(net917_c1,net917);
INTERCONNECT SplitCLK_2_407_SplitCLK_4_587(net918_c1,net918);
INTERCONNECT SplitCLK_2_407_SplitCLK_2_715(net919_c1,net919);
INTERCONNECT SplitCLK_0_406_SplitCLK_4_539(net920_c1,net920);
INTERCONNECT SplitCLK_0_406_SplitCLK_4_633(net921_c1,net921);
INTERCONNECT SplitCLK_6_405_SplitCLK_4_397(net922_c1,net922);
INTERCONNECT SplitCLK_6_405_SplitCLK_2_404(net923_c1,net923);
INTERCONNECT SplitCLK_2_404_SplitCLK_0_400(net924_c1,net924);
INTERCONNECT SplitCLK_2_404_SplitCLK_2_403(net925_c1,net925);
INTERCONNECT SplitCLK_2_403_SplitCLK_0_401(net926_c1,net926);
INTERCONNECT SplitCLK_2_403_SplitCLK_6_402(net927_c1,net927);
INTERCONNECT SplitCLK_6_402_SplitCLK_4_629(net928_c1,net928);
INTERCONNECT SplitCLK_6_402_SplitCLK_2_637(net929_c1,net929);
INTERCONNECT SplitCLK_0_401_SplitCLK_4_533(net930_c1,net930);
INTERCONNECT SplitCLK_0_401_SplitCLK_2_567(net931_c1,net931);
INTERCONNECT SplitCLK_0_400_SplitCLK_0_398(net932_c1,net932);
INTERCONNECT SplitCLK_0_400_SplitCLK_6_399(net933_c1,net933);
INTERCONNECT SplitCLK_6_399_SplitCLK_2_695(net934_c1,net934);
INTERCONNECT SplitCLK_6_399_SplitCLK_4_753(net935_c1,net935);
INTERCONNECT SplitCLK_0_398_SplitCLK_4_529(net936_c1,net936);
INTERCONNECT SplitCLK_0_398_SplitCLK_2_565(net937_c1,net937);
INTERCONNECT SplitCLK_4_397_SplitCLK_0_393(net938_c1,net938);
INTERCONNECT SplitCLK_4_397_SplitCLK_4_396(net939_c1,net939);
INTERCONNECT SplitCLK_4_396_SplitCLK_4_394(net940_c1,net940);
INTERCONNECT SplitCLK_4_396_SplitCLK_6_395(net941_c1,net941);
INTERCONNECT SplitCLK_6_395_SplitCLK_2_585(net942_c1,net942);
INTERCONNECT SplitCLK_6_395_SplitCLK_4_586(net943_c1,net943);
INTERCONNECT SplitCLK_4_394_SplitCLK_2_568(net944_c1,net944);
INTERCONNECT SplitCLK_4_394_SplitCLK_4_705(net945_c1,net945);
INTERCONNECT SplitCLK_0_393_SplitCLK_0_391(net946_c1,net946);
INTERCONNECT SplitCLK_0_393_SplitCLK_2_392(net947_c1,net947);
INTERCONNECT SplitCLK_2_392_SplitCLK_4_730(net948_c1,net948);
INTERCONNECT SplitCLK_2_392_SplitCLK_2_759(net949_c1,net949);
INTERCONNECT SplitCLK_0_391_SplitCLK_4_737(net950_c1,net950);
INTERCONNECT SplitCLK_0_391_SplitCLK_0_390(net951_c1,net951);
INTERCONNECT SplitCLK_0_390_DFFT_256__FPB_n715(net952_c1,net952);
INTERCONNECT SplitCLK_0_390_DFFT_257__FPB_n716(net953_c1,net953);
INTERCONNECT SplitCLK_0_389_SplitCLK_6_324(net954_c1,net954);
INTERCONNECT SplitCLK_0_389_SplitCLK_4_388(net955_c1,net955);
INTERCONNECT SplitCLK_4_388_SplitCLK_4_356(net956_c1,net956);
INTERCONNECT SplitCLK_4_388_SplitCLK_2_387(net957_c1,net957);
INTERCONNECT SplitCLK_2_387_SplitCLK_6_371(net958_c1,net958);
INTERCONNECT SplitCLK_2_387_SplitCLK_4_386(net959_c1,net959);
INTERCONNECT SplitCLK_4_386_SplitCLK_0_378(net960_c1,net960);
INTERCONNECT SplitCLK_4_386_SplitCLK_4_385(net961_c1,net961);
INTERCONNECT SplitCLK_4_385_SplitCLK_2_381(net962_c1,net962);
INTERCONNECT SplitCLK_4_385_SplitCLK_2_384(net963_c1,net963);
INTERCONNECT SplitCLK_2_384_SplitCLK_0_382(net964_c1,net964);
INTERCONNECT SplitCLK_2_384_SplitCLK_2_383(net965_c1,net965);
INTERCONNECT SplitCLK_2_383_SplitCLK_4_708(net966_c1,net966);
INTERCONNECT SplitCLK_2_383_SplitCLK_2_767(net967_c1,net967);
INTERCONNECT SplitCLK_0_382_SplitCLK_4_699(net968_c1,net968);
INTERCONNECT SplitCLK_0_382_SplitCLK_2_769(net969_c1,net969);
INTERCONNECT SplitCLK_2_381_SplitCLK_0_379(net970_c1,net970);
INTERCONNECT SplitCLK_2_381_SplitCLK_4_380(net971_c1,net971);
INTERCONNECT SplitCLK_4_380_SplitCLK_2_577(net972_c1,net972);
INTERCONNECT SplitCLK_4_380_SplitCLK_2_656(net973_c1,net973);
INTERCONNECT SplitCLK_0_379_SplitCLK_4_734(net974_c1,net974);
INTERCONNECT SplitCLK_0_379_SplitCLK_2_748(net975_c1,net975);
INTERCONNECT SplitCLK_0_378_SplitCLK_2_374(net976_c1,net976);
INTERCONNECT SplitCLK_0_378_SplitCLK_4_377(net977_c1,net977);
INTERCONNECT SplitCLK_4_377_SplitCLK_0_375(net978_c1,net978);
INTERCONNECT SplitCLK_4_377_SplitCLK_4_376(net979_c1,net979);
INTERCONNECT SplitCLK_4_376_SplitCLK_2_688(net980_c1,net980);
INTERCONNECT SplitCLK_4_376_SplitCLK_2_738(net981_c1,net981);
INTERCONNECT SplitCLK_0_375_SplitCLK_4_634(net982_c1,net982);
INTERCONNECT SplitCLK_0_375_SplitCLK_4_668(net983_c1,net983);
INTERCONNECT SplitCLK_2_374_SplitCLK_0_372(net984_c1,net984);
INTERCONNECT SplitCLK_2_374_SplitCLK_6_373(net985_c1,net985);
INTERCONNECT SplitCLK_6_373_SplitCLK_2_519(net986_c1,net986);
INTERCONNECT SplitCLK_6_373_SplitCLK_4_598(net987_c1,net987);
INTERCONNECT SplitCLK_0_372_SplitCLK_2_549(net988_c1,net988);
INTERCONNECT SplitCLK_0_372_SplitCLK_4_760(net989_c1,net989);
INTERCONNECT SplitCLK_6_371_SplitCLK_0_363(net990_c1,net990);
INTERCONNECT SplitCLK_6_371_SplitCLK_2_370(net991_c1,net991);
INTERCONNECT SplitCLK_2_370_SplitCLK_4_366(net992_c1,net992);
INTERCONNECT SplitCLK_2_370_SplitCLK_4_369(net993_c1,net993);
INTERCONNECT SplitCLK_4_369_SplitCLK_4_367(net994_c1,net994);
INTERCONNECT SplitCLK_4_369_SplitCLK_0_368(net995_c1,net995);
INTERCONNECT SplitCLK_0_368_SplitCLK_2_658(net996_c1,net996);
INTERCONNECT SplitCLK_0_368_SplitCLK_4_741(net997_c1,net997);
INTERCONNECT SplitCLK_4_367_SplitCLK_4_579(net998_c1,net998);
INTERCONNECT SplitCLK_4_367_SplitCLK_2_764(net999_c1,net999);
INTERCONNECT SplitCLK_4_366_SplitCLK_0_364(net1000_c1,net1000);
INTERCONNECT SplitCLK_4_366_SplitCLK_6_365(net1001_c1,net1001);
INTERCONNECT SplitCLK_6_365_SplitCLK_4_602(net1002_c1,net1002);
INTERCONNECT SplitCLK_6_365_SplitCLK_2_621(net1003_c1,net1003);
INTERCONNECT SplitCLK_0_364_SplitCLK_4_600(net1004_c1,net1004);
INTERCONNECT SplitCLK_0_364_SplitCLK_2_652(net1005_c1,net1005);
INTERCONNECT SplitCLK_0_363_SplitCLK_4_359(net1006_c1,net1006);
INTERCONNECT SplitCLK_0_363_SplitCLK_4_362(net1007_c1,net1007);
INTERCONNECT SplitCLK_4_362_SplitCLK_0_360(net1008_c1,net1008);
INTERCONNECT SplitCLK_4_362_SplitCLK_2_361(net1009_c1,net1009);
INTERCONNECT SplitCLK_2_361_SplitCLK_2_580(net1010_c1,net1010);
INTERCONNECT SplitCLK_2_361_SplitCLK_4_655(net1011_c1,net1011);
INTERCONNECT SplitCLK_0_360_SplitCLK_4_662(net1012_c1,net1012);
INTERCONNECT SplitCLK_0_360_SplitCLK_2_696(net1013_c1,net1013);
INTERCONNECT SplitCLK_4_359_SplitCLK_0_357(net1014_c1,net1014);
INTERCONNECT SplitCLK_4_359_SplitCLK_6_358(net1015_c1,net1015);
INTERCONNECT SplitCLK_6_358_SplitCLK_4_603(net1016_c1,net1016);
INTERCONNECT SplitCLK_6_358_SplitCLK_2_635(net1017_c1,net1017);
INTERCONNECT SplitCLK_0_357_SplitCLK_2_657(net1018_c1,net1018);
INTERCONNECT SplitCLK_0_357_SplitCLK_4_678(net1019_c1,net1019);
INTERCONNECT SplitCLK_4_356_SplitCLK_6_340(net1020_c1,net1020);
INTERCONNECT SplitCLK_4_356_SplitCLK_4_355(net1021_c1,net1021);
INTERCONNECT SplitCLK_4_355_SplitCLK_0_347(net1022_c1,net1022);
INTERCONNECT SplitCLK_4_355_SplitCLK_4_354(net1023_c1,net1023);
INTERCONNECT SplitCLK_4_354_SplitCLK_6_350(net1024_c1,net1024);
INTERCONNECT SplitCLK_4_354_SplitCLK_4_353(net1025_c1,net1025);
INTERCONNECT SplitCLK_4_353_SplitCLK_4_351(net1026_c1,net1026);
INTERCONNECT SplitCLK_4_353_SplitCLK_2_352(net1027_c1,net1027);
INTERCONNECT SplitCLK_2_352_SplitCLK_4_589(net1028_c1,net1028);
INTERCONNECT SplitCLK_2_352_SplitCLK_2_754(net1029_c1,net1029);
INTERCONNECT SplitCLK_4_351_SplitCLK_2_666(net1030_c1,net1030);
INTERCONNECT SplitCLK_4_351_SplitCLK_4_686(net1031_c1,net1031);
INTERCONNECT SplitCLK_6_350_SplitCLK_0_348(net1032_c1,net1032);
INTERCONNECT SplitCLK_6_350_SplitCLK_6_349(net1033_c1,net1033);
INTERCONNECT SplitCLK_6_349_SplitCLK_4_762(net1034_c1,net1034);
INTERCONNECT SplitCLK_6_349_SplitCLK_2_763(net1035_c1,net1035);
INTERCONNECT SplitCLK_0_348_SplitCLK_4_750(net1036_c1,net1036);
INTERCONNECT SplitCLK_0_348_SplitCLK_4_756(net1037_c1,net1037);
INTERCONNECT SplitCLK_0_347_SplitCLK_4_343(net1038_c1,net1038);
INTERCONNECT SplitCLK_0_347_SplitCLK_4_346(net1039_c1,net1039);
INTERCONNECT SplitCLK_4_346_SplitCLK_0_344(net1040_c1,net1040);
INTERCONNECT SplitCLK_4_346_SplitCLK_4_345(net1041_c1,net1041);
INTERCONNECT SplitCLK_4_345_SplitCLK_2_697(net1042_c1,net1042);
INTERCONNECT SplitCLK_4_345_SplitCLK_2_727(net1043_c1,net1043);
INTERCONNECT SplitCLK_0_344_SplitCLK_4_706(net1044_c1,net1044);
INTERCONNECT SplitCLK_0_344_SplitCLK_4_718(net1045_c1,net1045);
INTERCONNECT SplitCLK_4_343_SplitCLK_4_341(net1046_c1,net1046);
INTERCONNECT SplitCLK_4_343_SplitCLK_6_342(net1047_c1,net1047);
INTERCONNECT SplitCLK_6_342_SplitCLK_2_665(net1048_c1,net1048);
INTERCONNECT SplitCLK_6_342_SplitCLK_4_683(net1049_c1,net1049);
INTERCONNECT SplitCLK_4_341_SplitCLK_2_692(net1050_c1,net1050);
INTERCONNECT SplitCLK_4_341_SplitCLK_4_703(net1051_c1,net1051);
INTERCONNECT SplitCLK_6_340_SplitCLK_4_332(net1052_c1,net1052);
INTERCONNECT SplitCLK_6_340_SplitCLK_6_339(net1053_c1,net1053);
INTERCONNECT SplitCLK_6_339_SplitCLK_6_335(net1054_c1,net1054);
INTERCONNECT SplitCLK_6_339_SplitCLK_4_338(net1055_c1,net1055);
INTERCONNECT SplitCLK_4_338_SplitCLK_4_336(net1056_c1,net1056);
INTERCONNECT SplitCLK_4_338_SplitCLK_2_337(net1057_c1,net1057);
INTERCONNECT SplitCLK_2_337_SplitCLK_4_559(net1058_c1,net1058);
INTERCONNECT SplitCLK_2_337_SplitCLK_2_661(net1059_c1,net1059);
INTERCONNECT SplitCLK_4_336_SplitCLK_2_581(net1060_c1,net1060);
INTERCONNECT SplitCLK_4_336_SplitCLK_4_583(net1061_c1,net1061);
INTERCONNECT SplitCLK_6_335_SplitCLK_0_333(net1062_c1,net1062);
INTERCONNECT SplitCLK_6_335_SplitCLK_6_334(net1063_c1,net1063);
INTERCONNECT SplitCLK_6_334_SplitCLK_2_575(net1064_c1,net1064);
INTERCONNECT SplitCLK_6_334_SplitCLK_4_660(net1065_c1,net1065);
INTERCONNECT SplitCLK_0_333_SplitCLK_4_676(net1066_c1,net1066);
INTERCONNECT SplitCLK_0_333_SplitCLK_4_768(net1067_c1,net1067);
INTERCONNECT SplitCLK_4_332_SplitCLK_0_328(net1068_c1,net1068);
INTERCONNECT SplitCLK_4_332_SplitCLK_4_331(net1069_c1,net1069);
INTERCONNECT SplitCLK_4_331_SplitCLK_0_329(net1070_c1,net1070);
INTERCONNECT SplitCLK_4_331_SplitCLK_2_330(net1071_c1,net1071);
INTERCONNECT SplitCLK_2_330_SplitCLK_2_582(net1072_c1,net1072);
INTERCONNECT SplitCLK_2_330_SplitCLK_4_765(net1073_c1,net1073);
INTERCONNECT SplitCLK_0_329_SplitCLK_4_546(net1074_c1,net1074);
INTERCONNECT SplitCLK_0_329_SplitCLK_2_571(net1075_c1,net1075);
INTERCONNECT SplitCLK_0_328_SplitCLK_2_326(net1076_c1,net1076);
INTERCONNECT SplitCLK_0_328_SplitCLK_6_327(net1077_c1,net1077);
INTERCONNECT SplitCLK_6_327_SplitCLK_2_672(net1078_c1,net1078);
INTERCONNECT SplitCLK_6_327_SplitCLK_2_713(net1079_c1,net1079);
INTERCONNECT SplitCLK_2_326_SplitCLK_2_560(net1080_c1,net1080);
INTERCONNECT SplitCLK_2_326_SplitCLK_4_325(net1081_c1,net1081);
INTERCONNECT SplitCLK_4_325_AND2T_38_n74(net1082_c1,net1082);
INTERCONNECT SplitCLK_4_325_DFFT_166__FPB_n625(net1083_c1,net1083);
INTERCONNECT SplitCLK_6_324_SplitCLK_0_292(net1084_c1,net1084);
INTERCONNECT SplitCLK_6_324_SplitCLK_2_323(net1085_c1,net1085);
INTERCONNECT SplitCLK_2_323_SplitCLK_2_307(net1086_c1,net1086);
INTERCONNECT SplitCLK_2_323_SplitCLK_4_322(net1087_c1,net1087);
INTERCONNECT SplitCLK_4_322_SplitCLK_0_314(net1088_c1,net1088);
INTERCONNECT SplitCLK_4_322_SplitCLK_2_321(net1089_c1,net1089);
INTERCONNECT SplitCLK_2_321_SplitCLK_6_317(net1090_c1,net1090);
INTERCONNECT SplitCLK_2_321_SplitCLK_4_320(net1091_c1,net1091);
INTERCONNECT SplitCLK_4_320_SplitCLK_4_318(net1092_c1,net1092);
INTERCONNECT SplitCLK_4_320_SplitCLK_2_319(net1093_c1,net1093);
INTERCONNECT SplitCLK_2_319_SplitCLK_4_547(net1094_c1,net1094);
INTERCONNECT SplitCLK_2_319_SplitCLK_2_702(net1095_c1,net1095);
INTERCONNECT SplitCLK_4_318_SplitCLK_2_563(net1096_c1,net1096);
INTERCONNECT SplitCLK_4_318_SplitCLK_4_651(net1097_c1,net1097);
INTERCONNECT SplitCLK_6_317_SplitCLK_4_315(net1098_c1,net1098);
INTERCONNECT SplitCLK_6_317_SplitCLK_6_316(net1099_c1,net1099);
INTERCONNECT SplitCLK_6_316_SplitCLK_2_537(net1100_c1,net1100);
INTERCONNECT SplitCLK_6_316_SplitCLK_2_553(net1101_c1,net1101);
INTERCONNECT SplitCLK_4_315_SplitCLK_2_525(net1102_c1,net1102);
INTERCONNECT SplitCLK_4_315_SplitCLK_2_526(net1103_c1,net1103);
INTERCONNECT SplitCLK_0_314_SplitCLK_6_310(net1104_c1,net1104);
INTERCONNECT SplitCLK_0_314_SplitCLK_4_313(net1105_c1,net1105);
INTERCONNECT SplitCLK_4_313_SplitCLK_4_311(net1106_c1,net1106);
INTERCONNECT SplitCLK_4_313_SplitCLK_6_312(net1107_c1,net1107);
INTERCONNECT SplitCLK_6_312_SplitCLK_4_574(net1108_c1,net1108);
INTERCONNECT SplitCLK_6_312_SplitCLK_2_757(net1109_c1,net1109);
INTERCONNECT SplitCLK_4_311_SplitCLK_4_561(net1110_c1,net1110);
INTERCONNECT SplitCLK_4_311_SplitCLK_4_578(net1111_c1,net1111);
INTERCONNECT SplitCLK_6_310_SplitCLK_0_308(net1112_c1,net1112);
INTERCONNECT SplitCLK_6_310_SplitCLK_6_309(net1113_c1,net1113);
INTERCONNECT SplitCLK_6_309_SplitCLK_4_588(net1114_c1,net1114);
INTERCONNECT SplitCLK_6_309_SplitCLK_2_654(net1115_c1,net1115);
INTERCONNECT SplitCLK_0_308_SplitCLK_4_726(net1116_c1,net1116);
INTERCONNECT SplitCLK_0_308_SplitCLK_4_735(net1117_c1,net1117);
INTERCONNECT SplitCLK_2_307_SplitCLK_4_299(net1118_c1,net1118);
INTERCONNECT SplitCLK_2_307_SplitCLK_6_306(net1119_c1,net1119);
INTERCONNECT SplitCLK_6_306_SplitCLK_2_302(net1120_c1,net1120);
INTERCONNECT SplitCLK_6_306_SplitCLK_4_305(net1121_c1,net1121);
INTERCONNECT SplitCLK_4_305_SplitCLK_0_303(net1122_c1,net1122);
INTERCONNECT SplitCLK_4_305_SplitCLK_2_304(net1123_c1,net1123);
INTERCONNECT SplitCLK_2_304_SplitCLK_4_532(net1124_c1,net1124);
INTERCONNECT SplitCLK_2_304_SplitCLK_2_747(net1125_c1,net1125);
INTERCONNECT SplitCLK_0_303_SplitCLK_2_530(net1126_c1,net1126);
INTERCONNECT SplitCLK_0_303_SplitCLK_4_700(net1127_c1,net1127);
INTERCONNECT SplitCLK_2_302_SplitCLK_0_300(net1128_c1,net1128);
INTERCONNECT SplitCLK_2_302_SplitCLK_6_301(net1129_c1,net1129);
INTERCONNECT SplitCLK_6_301_SplitCLK_2_566(net1130_c1,net1130);
INTERCONNECT SplitCLK_6_301_SplitCLK_4_758(net1131_c1,net1131);
INTERCONNECT SplitCLK_0_300_SplitCLK_4_594(net1132_c1,net1132);
INTERCONNECT SplitCLK_0_300_SplitCLK_2_752(net1133_c1,net1133);
INTERCONNECT SplitCLK_4_299_SplitCLK_6_295(net1134_c1,net1134);
INTERCONNECT SplitCLK_4_299_SplitCLK_0_298(net1135_c1,net1135);
INTERCONNECT SplitCLK_0_298_SplitCLK_4_296(net1136_c1,net1136);
INTERCONNECT SplitCLK_0_298_SplitCLK_4_297(net1137_c1,net1137);
INTERCONNECT SplitCLK_4_297_SplitCLK_2_570(net1138_c1,net1138);
INTERCONNECT SplitCLK_4_297_SplitCLK_2_648(net1139_c1,net1139);
INTERCONNECT SplitCLK_4_296_SplitCLK_2_542(net1140_c1,net1140);
INTERCONNECT SplitCLK_4_296_SplitCLK_4_544(net1141_c1,net1141);
INTERCONNECT SplitCLK_6_295_SplitCLK_4_293(net1142_c1,net1142);
INTERCONNECT SplitCLK_6_295_SplitCLK_6_294(net1143_c1,net1143);
INTERCONNECT SplitCLK_6_294_SplitCLK_4_710(net1144_c1,net1144);
INTERCONNECT SplitCLK_6_294_SplitCLK_2_746(net1145_c1,net1145);
INTERCONNECT SplitCLK_4_293_SplitCLK_2_721(net1146_c1,net1146);
INTERCONNECT SplitCLK_4_293_SplitCLK_4_729(net1147_c1,net1147);
INTERCONNECT SplitCLK_0_292_SplitCLK_6_276(net1148_c1,net1148);
INTERCONNECT SplitCLK_0_292_SplitCLK_4_291(net1149_c1,net1149);
INTERCONNECT SplitCLK_4_291_SplitCLK_0_283(net1150_c1,net1150);
INTERCONNECT SplitCLK_4_291_SplitCLK_2_290(net1151_c1,net1151);
INTERCONNECT SplitCLK_2_290_SplitCLK_6_286(net1152_c1,net1152);
INTERCONNECT SplitCLK_2_290_SplitCLK_4_289(net1153_c1,net1153);
INTERCONNECT SplitCLK_4_289_SplitCLK_0_287(net1154_c1,net1154);
INTERCONNECT SplitCLK_4_289_SplitCLK_2_288(net1155_c1,net1155);
INTERCONNECT SplitCLK_2_288_SplitCLK_2_551(net1156_c1,net1156);
INTERCONNECT SplitCLK_2_288_SplitCLK_2_562(net1157_c1,net1157);
INTERCONNECT SplitCLK_0_287_SplitCLK_4_543(net1158_c1,net1158);
INTERCONNECT SplitCLK_0_287_SplitCLK_4_557(net1159_c1,net1159);
INTERCONNECT SplitCLK_6_286_SplitCLK_0_284(net1160_c1,net1160);
INTERCONNECT SplitCLK_6_286_SplitCLK_4_285(net1161_c1,net1161);
INTERCONNECT SplitCLK_4_285_SplitCLK_2_524(net1162_c1,net1162);
INTERCONNECT SplitCLK_4_285_SplitCLK_2_714(net1163_c1,net1163);
INTERCONNECT SplitCLK_0_284_SplitCLK_4_639(net1164_c1,net1164);
INTERCONNECT SplitCLK_0_284_SplitCLK_4_693(net1165_c1,net1165);
INTERCONNECT SplitCLK_0_283_SplitCLK_4_279(net1166_c1,net1166);
INTERCONNECT SplitCLK_0_283_SplitCLK_4_282(net1167_c1,net1167);
INTERCONNECT SplitCLK_4_282_SplitCLK_0_280(net1168_c1,net1168);
INTERCONNECT SplitCLK_4_282_SplitCLK_0_281(net1169_c1,net1169);
INTERCONNECT SplitCLK_0_281_SplitCLK_4_555(net1170_c1,net1170);
INTERCONNECT SplitCLK_0_281_SplitCLK_4_576(net1171_c1,net1171);
INTERCONNECT SplitCLK_0_280_SplitCLK_2_550(net1172_c1,net1172);
INTERCONNECT SplitCLK_0_280_SplitCLK_4_552(net1173_c1,net1173);
INTERCONNECT SplitCLK_4_279_SplitCLK_0_277(net1174_c1,net1174);
INTERCONNECT SplitCLK_4_279_SplitCLK_2_278(net1175_c1,net1175);
INTERCONNECT SplitCLK_2_278_SplitCLK_2_569(net1176_c1,net1176);
INTERCONNECT SplitCLK_2_278_SplitCLK_2_638(net1177_c1,net1177);
INTERCONNECT SplitCLK_0_277_SplitCLK_4_724(net1178_c1,net1178);
INTERCONNECT SplitCLK_0_277_SplitCLK_2_743(net1179_c1,net1179);
INTERCONNECT SplitCLK_6_276_SplitCLK_4_268(net1180_c1,net1180);
INTERCONNECT SplitCLK_6_276_SplitCLK_2_275(net1181_c1,net1181);
INTERCONNECT SplitCLK_2_275_SplitCLK_6_271(net1182_c1,net1182);
INTERCONNECT SplitCLK_2_275_SplitCLK_4_274(net1183_c1,net1183);
INTERCONNECT SplitCLK_4_274_SplitCLK_0_272(net1184_c1,net1184);
INTERCONNECT SplitCLK_4_274_SplitCLK_2_273(net1185_c1,net1185);
INTERCONNECT SplitCLK_2_273_SplitCLK_2_591(net1186_c1,net1186);
INTERCONNECT SplitCLK_2_273_SplitCLK_2_709(net1187_c1,net1187);
INTERCONNECT SplitCLK_0_272_SplitCLK_2_663(net1188_c1,net1188);
INTERCONNECT SplitCLK_0_272_SplitCLK_4_704(net1189_c1,net1189);
INTERCONNECT SplitCLK_6_271_SplitCLK_0_269(net1190_c1,net1190);
INTERCONNECT SplitCLK_6_271_SplitCLK_6_270(net1191_c1,net1191);
INTERCONNECT SplitCLK_6_270_SplitCLK_4_595(net1192_c1,net1192);
INTERCONNECT SplitCLK_6_270_SplitCLK_2_736(net1193_c1,net1193);
INTERCONNECT SplitCLK_0_269_SplitCLK_2_531(net1194_c1,net1194);
INTERCONNECT SplitCLK_0_269_SplitCLK_4_647(net1195_c1,net1195);
INTERCONNECT SplitCLK_4_268_SplitCLK_0_264(net1196_c1,net1196);
INTERCONNECT SplitCLK_4_268_SplitCLK_6_267(net1197_c1,net1197);
INTERCONNECT SplitCLK_6_267_SplitCLK_0_265(net1198_c1,net1198);
INTERCONNECT SplitCLK_6_267_SplitCLK_2_266(net1199_c1,net1199);
INTERCONNECT SplitCLK_2_266_SplitCLK_4_534(net1200_c1,net1200);
INTERCONNECT SplitCLK_2_266_SplitCLK_2_640(net1201_c1,net1201);
INTERCONNECT SplitCLK_0_265_SplitCLK_4_527(net1202_c1,net1202);
INTERCONNECT SplitCLK_0_265_SplitCLK_4_617(net1203_c1,net1203);
INTERCONNECT SplitCLK_0_264_SplitCLK_0_262(net1204_c1,net1204);
INTERCONNECT SplitCLK_0_264_SplitCLK_6_263(net1205_c1,net1205);
INTERCONNECT SplitCLK_6_263_SplitCLK_2_716(net1206_c1,net1206);
INTERCONNECT SplitCLK_6_263_SplitCLK_4_720(net1207_c1,net1207);
INTERCONNECT SplitCLK_0_262_SplitCLK_4_631(net1208_c1,net1208);
INTERCONNECT SplitCLK_0_262_SplitCLK_0_261(net1209_c1,net1209);
INTERCONNECT SplitCLK_0_261_DFFT_262__FPB_n721(net1210_c1,net1210);
INTERCONNECT SplitCLK_0_261_DFFT_263__FPB_n722(net1211_c1,net1211);
INTERCONNECT GCLK_Pad_SplitCLK_0_771(GCLK_Pad,net1212);
INTERCONNECT Split_HOLD_869_DFFT_189__FPB_n648(net1213_c1,net1213);
INTERCONNECT Split_HOLD_870_DFFT_237__FPB_n696(net1214_c1,net1214);
INTERCONNECT Split_HOLD_871_OR2T_80_n116(net1215_c1,net1215);
INTERCONNECT Split_HOLD_872_DFFT_152__FPB_n611(net1216_c1,net1216);
INTERCONNECT Split_HOLD_873_DFFT_223__FPB_n682(net1217_c1,net1217);
INTERCONNECT Split_HOLD_874_DFFT_201__FPB_n660(net1218_c1,net1218);
INTERCONNECT Split_HOLD_875_AND2T_67_n103(net1219_c1,net1219);
INTERCONNECT Split_HOLD_876_AND2T_92_n128(net1220_c1,net1220);
INTERCONNECT Split_HOLD_877_AND2T_49_n85(net1221_c1,net1221);

endmodule
