module counter1_route(
input GCLK_Pad,
input en_Pad,
input rst_Pad,
output count_Pad);

wire net0_c1;
wire net0;
wire net1_c1;
wire net1;
wire en_Pad;
wire net2;
wire net3_c1;
wire net3;
wire rst_Pad;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire count_Pad;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire GCLK_Pad;
wire net14;

AND2T AND2T_7_n10(net10,net1,net0,net3_c1);
XOR2T XOR2T_6_n9(net12,net5,net2,net1_c1);
DFFT DFFT_8__FBL_n11(net13,net3,net7_c1);
NOTT NOTT_5_n8(net11,net4,net0_c1);
SPLITT Split_9_count(net7,net5_c1,net6_c1);
SPLITT SplitCLK_4_5(net8,net12_c1,net13_c1);
SPLITT SplitCLK_4_6(net9,net10_c1,net11_c1);
SPLITT SplitCLK_0_7(net14,net8_c1,net9_c1);
INTERCONNECT NOTT_5_n8_AND2T_7_n10(net0_c1,net0);
INTERCONNECT XOR2T_6_n9_AND2T_7_n10(net1_c1,net1);
INTERCONNECT en_Pad_XOR2T_6_n9(en_Pad,net2);
INTERCONNECT AND2T_7_n10_DFFT_8__FBL_n11(net3_c1,net3);
INTERCONNECT rst_Pad_NOTT_5_n8(rst_Pad,net4);
INTERCONNECT Split_9_count_XOR2T_6_n9(net5_c1,net5);
INTERCONNECT Split_9_count_count_Pad(net6_c1,count_Pad);
INTERCONNECT DFFT_8__FBL_n11_Split_9_count(net7_c1,net7);
INTERCONNECT SplitCLK_0_7_SplitCLK_4_5(net8_c1,net8);
INTERCONNECT SplitCLK_0_7_SplitCLK_4_6(net9_c1,net9);
INTERCONNECT SplitCLK_4_6_AND2T_7_n10(net10_c1,net10);
INTERCONNECT SplitCLK_4_6_NOTT_5_n8(net11_c1,net11);
INTERCONNECT SplitCLK_4_5_XOR2T_6_n9(net12_c1,net12);
INTERCONNECT SplitCLK_4_5_DFFT_8__FBL_n11(net13_c1,net13);
INTERCONNECT GCLK_Pad_SplitCLK_0_7(GCLK_Pad,net14);

endmodule
