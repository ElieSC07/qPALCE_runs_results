module TAP_route(
input GCLK_Pad,
input TMS_Pad,
output TDO_Pad);

wire net0_c1;
wire net0;
wire TMS_Pad;
wire net1;
wire net2_c1;
wire net2;
wire net3_c1;
wire net3;
wire net4_c1;
wire net4;
wire net5_c1;
wire net5;
wire net6_c1;
wire net6;
wire net7_c1;
wire net7;
wire net8_c1;
wire net8;
wire net9_c1;
wire net9;
wire net10_c1;
wire net10;
wire net11_c1;
wire net11;
wire net12_c1;
wire net12;
wire net13_c1;
wire net13;
wire net14_c1;
wire net14;
wire net15_c1;
wire net15;
wire net16_c1;
wire net16;
wire net17_c1;
wire net17;
wire net18_c1;
wire net18;
wire net19_c1;
wire net19;
wire net20_c1;
wire net20;
wire net21_c1;
wire net21;
wire net22_c1;
wire net22;
wire net23_c1;
wire net23;
wire net24_c1;
wire net24;
wire net25_c1;
wire net25;
wire net26_c1;
wire net26;
wire net27_c1;
wire net27;
wire net28_c1;
wire net28;
wire net29_c1;
wire net29;
wire net30_c1;
wire net30;
wire net31_c1;
wire net31;
wire net32_c1;
wire net32;
wire net33_c1;
wire net33;
wire net34_c1;
wire net34;
wire net35_c1;
wire net35;
wire net36_c1;
wire net36;
wire net37_c1;
wire net37;
wire net38_c1;
wire net38;
wire net39_c1;
wire net39;
wire net40_c1;
wire net40;
wire net41_c1;
wire net41;
wire net42_c1;
wire net42;
wire net43_c1;
wire net43;
wire net44_c1;
wire net44;
wire net45_c1;
wire net45;
wire net46_c1;
wire net46;
wire net47_c1;
wire net47;
wire net48_c1;
wire net48;
wire net49_c1;
wire net49;
wire net50_c1;
wire net50;
wire net51_c1;
wire net51;
wire net52_c1;
wire net52;
wire net53_c1;
wire net53;
wire net54_c1;
wire net54;
wire net55_c1;
wire net55;
wire net56_c1;
wire net56;
wire net57_c1;
wire net57;
wire net58_c1;
wire net58;
wire net59_c1;
wire net59;
wire net60_c1;
wire net60;
wire net61_c1;
wire net61;
wire net62_c1;
wire net62;
wire net63_c1;
wire net63;
wire net64_c1;
wire net64;
wire net65_c1;
wire net65;
wire net66_c1;
wire net66;
wire net67_c1;
wire net67;
wire net68_c1;
wire net68;
wire net69_c1;
wire net69;
wire net70_c1;
wire net70;
wire net71_c1;
wire net71;
wire net72_c1;
wire net72;
wire net73_c1;
wire net73;
wire net74_c1;
wire net74;
wire net75_c1;
wire net75;
wire net76_c1;
wire net76;
wire net77_c1;
wire net77;
wire net78_c1;
wire net78;
wire net79_c1;
wire net79;
wire net80_c1;
wire net80;
wire net81_c1;
wire net81;
wire net82_c1;
wire net82;
wire net83_c1;
wire net83;
wire net84_c1;
wire net84;
wire net85_c1;
wire net85;
wire net86_c1;
wire net86;
wire net87_c1;
wire net87;
wire net88_c1;
wire net88;
wire net89_c1;
wire net89;
wire net90_c1;
wire net90;
wire net91_c1;
wire net91;
wire net92_c1;
wire net92;
wire net93_c1;
wire net93;
wire net94_c1;
wire net94;
wire net95_c1;
wire net95;
wire net96_c1;
wire net96;
wire net97_c1;
wire net97;
wire net98_c1;
wire net98;
wire net99_c1;
wire net99;
wire net100_c1;
wire net100;
wire net101_c1;
wire net101;
wire net102_c1;
wire net102;
wire net103_c1;
wire net103;
wire net104_c1;
wire net104;
wire net105_c1;
wire net105;
wire net106_c1;
wire net106;
wire net107_c1;
wire net107;
wire net108_c1;
wire net108;
wire net109_c1;
wire net109;
wire net110_c1;
wire net110;
wire net111_c1;
wire net111;
wire net112_c1;
wire net112;
wire net113_c1;
wire net113;
wire net114_c1;
wire net114;
wire net115_c1;
wire net115;
wire net116_c1;
wire net116;
wire net117_c1;
wire net117;
wire net118_c1;
wire net118;
wire net119_c1;
wire net119;
wire net120_c1;
wire net120;
wire net121_c1;
wire net121;
wire net122_c1;
wire net122;
wire net123_c1;
wire net123;
wire net124_c1;
wire net124;
wire net125_c1;
wire net125;
wire net126_c1;
wire net126;
wire net127_c1;
wire net127;
wire net128_c1;
wire net128;
wire net129_c1;
wire net129;
wire net130_c1;
wire net130;
wire net131_c1;
wire net131;
wire net132_c1;
wire net132;
wire net133_c1;
wire net133;
wire net134_c1;
wire net134;
wire net135_c1;
wire net135;
wire net136_c1;
wire net136;
wire net137_c1;
wire net137;
wire net138_c1;
wire net138;
wire net139_c1;
wire net139;
wire net140_c1;
wire net140;
wire net141_c1;
wire net141;
wire net142_c1;
wire net142;
wire net143_c1;
wire net143;
wire net144_c1;
wire net144;
wire net145_c1;
wire net145;
wire net146_c1;
wire net146;
wire net147_c1;
wire net147;
wire net148_c1;
wire net148;
wire net149_c1;
wire net149;
wire net150_c1;
wire net150;
wire net151_c1;
wire net151;
wire net152_c1;
wire net152;
wire net153_c1;
wire net153;
wire net154_c1;
wire net154;
wire net155_c1;
wire net155;
wire net156_c1;
wire net156;
wire net157_c1;
wire net157;
wire net158_c1;
wire net158;
wire net159_c1;
wire net159;
wire net160_c1;
wire net160;
wire net161_c1;
wire net161;
wire net162_c1;
wire net162;
wire net163_c1;
wire net163;
wire net164_c1;
wire net164;
wire net165_c1;
wire net165;
wire net166_c1;
wire net166;
wire net167_c1;
wire net167;
wire net168_c1;
wire net168;
wire net169_c1;
wire net169;
wire net170_c1;
wire net170;
wire net171_c1;
wire net171;
wire net172_c1;
wire net172;
wire net173_c1;
wire net173;
wire net174_c1;
wire net174;
wire net175_c1;
wire net175;
wire net176_c1;
wire net176;
wire net177_c1;
wire net177;
wire net178_c1;
wire net178;
wire net179_c1;
wire net179;
wire net180_c1;
wire net180;
wire net181_c1;
wire net181;
wire net182_c1;
wire net182;
wire net183_c1;
wire net183;
wire net184_c1;
wire net184;
wire net185_c1;
wire net185;
wire net186_c1;
wire net186;
wire net187_c1;
wire net187;
wire net188_c1;
wire net188;
wire net189_c1;
wire net189;
wire net190_c1;
wire net190;
wire net191_c1;
wire net191;
wire net192_c1;
wire net192;
wire net193_c1;
wire net193;
wire net194_c1;
wire net194;
wire net195_c1;
wire net195;
wire net196_c1;
wire net196;
wire net197_c1;
wire net197;
wire net198_c1;
wire net198;
wire net199_c1;
wire net199;
wire net200_c1;
wire net200;
wire net201_c1;
wire net201;
wire net202_c1;
wire net202;
wire net203_c1;
wire net203;
wire net204_c1;
wire net204;
wire net205_c1;
wire net205;
wire net206_c1;
wire net206;
wire net207_c1;
wire net207;
wire net208_c1;
wire net208;
wire net209_c1;
wire net209;
wire net210_c1;
wire net210;
wire net211_c1;
wire net211;
wire net212_c1;
wire net212;
wire net213_c1;
wire net213;
wire net214_c1;
wire net214;
wire net215_c1;
wire net215;
wire net216_c1;
wire net216;
wire net217_c1;
wire net217;
wire net218_c1;
wire net218;
wire net219_c1;
wire net219;
wire net220_c1;
wire net220;
wire net221_c1;
wire net221;
wire net222_c1;
wire net222;
wire net223_c1;
wire net223;
wire net224_c1;
wire net224;
wire net225_c1;
wire net225;
wire net226_c1;
wire net226;
wire net227_c1;
wire net227;
wire net228_c1;
wire net228;
wire net229_c1;
wire net229;
wire net230_c1;
wire net230;
wire net231_c1;
wire net231;
wire net232_c1;
wire net232;
wire net233_c1;
wire net233;
wire net234_c1;
wire net234;
wire net235_c1;
wire net235;
wire net236_c1;
wire net236;
wire net237_c1;
wire net237;
wire net238_c1;
wire net238;
wire net239_c1;
wire net239;
wire net240_c1;
wire net240;
wire net241_c1;
wire net241;
wire net242_c1;
wire net242;
wire net243_c1;
wire net243;
wire net244_c1;
wire net244;
wire net245_c1;
wire net245;
wire net246_c1;
wire net246;
wire net247_c1;
wire net247;
wire net248_c1;
wire net248;
wire net249_c1;
wire net249;
wire net250_c1;
wire net250;
wire net251_c1;
wire net251;
wire net252_c1;
wire net252;
wire net253_c1;
wire net253;
wire net254_c1;
wire net254;
wire net255_c1;
wire net255;
wire net256_c1;
wire net256;
wire net257_c1;
wire net257;
wire net258_c1;
wire net258;
wire net259_c1;
wire net259;
wire net260_c1;
wire net260;
wire net261_c1;
wire net261;
wire net262_c1;
wire net262;
wire net263_c1;
wire net263;
wire net264_c1;
wire net264;
wire net265_c1;
wire net265;
wire net266_c1;
wire TDO_Pad;
wire net267_c1;
wire net267;
wire net268_c1;
wire net268;
wire net269_c1;
wire net269;
wire net270_c1;
wire net270;
wire net271_c1;
wire net271;
wire net272_c1;
wire net272;
wire net273_c1;
wire net273;
wire net274_c1;
wire net274;
wire net275_c1;
wire net275;
wire net276_c1;
wire net276;
wire net277_c1;
wire net277;
wire net278_c1;
wire net278;
wire net279_c1;
wire net279;
wire net280_c1;
wire net280;
wire net281_c1;
wire net281;
wire net282_c1;
wire net282;
wire net283_c1;
wire net283;
wire net284_c1;
wire net284;
wire net285_c1;
wire net285;
wire net286_c1;
wire net286;
wire net287_c1;
wire net287;
wire net288_c1;
wire net288;
wire net289_c1;
wire net289;
wire net290_c1;
wire net290;
wire net291_c1;
wire net291;
wire net292_c1;
wire net292;
wire net293_c1;
wire net293;
wire net294_c1;
wire net294;
wire net295_c1;
wire net295;
wire net296_c1;
wire net296;
wire net297_c1;
wire net297;
wire net298_c1;
wire net298;
wire net299_c1;
wire net299;
wire net300_c1;
wire net300;
wire net301_c1;
wire net301;
wire net302_c1;
wire net302;
wire net303_c1;
wire net303;
wire net304_c1;
wire net304;
wire net305_c1;
wire net305;
wire net306_c1;
wire net306;
wire net307_c1;
wire net307;
wire net308_c1;
wire net308;
wire net309_c1;
wire net309;
wire net310_c1;
wire net310;
wire net311_c1;
wire net311;
wire net312_c1;
wire net312;
wire net313_c1;
wire net313;
wire net314_c1;
wire net314;
wire net315_c1;
wire net315;
wire net316_c1;
wire net316;
wire net317_c1;
wire net317;
wire net318_c1;
wire net318;
wire net319_c1;
wire net319;
wire net320_c1;
wire net320;
wire net321_c1;
wire net321;
wire net322_c1;
wire net322;
wire net323_c1;
wire net323;
wire net324_c1;
wire net324;
wire net325_c1;
wire net325;
wire net326_c1;
wire net326;
wire net327_c1;
wire net327;
wire net328_c1;
wire net328;
wire net329_c1;
wire net329;
wire net330_c1;
wire net330;
wire net331_c1;
wire net331;
wire net332_c1;
wire net332;
wire net333_c1;
wire net333;
wire net334_c1;
wire net334;
wire net335_c1;
wire net335;
wire net336_c1;
wire net336;
wire net337_c1;
wire net337;
wire net338_c1;
wire net338;
wire net339_c1;
wire net339;
wire net340_c1;
wire net340;
wire net341_c1;
wire net341;
wire net342_c1;
wire net342;
wire net343_c1;
wire net343;
wire net344_c1;
wire net344;
wire net345_c1;
wire net345;
wire net346_c1;
wire net346;
wire net347_c1;
wire net347;
wire net348_c1;
wire net348;
wire net349_c1;
wire net349;
wire net350_c1;
wire net350;
wire net351_c1;
wire net351;
wire net352_c1;
wire net352;
wire net353_c1;
wire net353;
wire net354_c1;
wire net354;
wire net355_c1;
wire net355;
wire net356_c1;
wire net356;
wire net357_c1;
wire net357;
wire net358_c1;
wire net358;
wire net359_c1;
wire net359;
wire net360_c1;
wire net360;
wire net361_c1;
wire net361;
wire net362_c1;
wire net362;
wire net363_c1;
wire net363;
wire net364_c1;
wire net364;
wire net365_c1;
wire net365;
wire net366_c1;
wire net366;
wire net367_c1;
wire net367;
wire net368_c1;
wire net368;
wire net369_c1;
wire net369;
wire net370_c1;
wire net370;
wire net371_c1;
wire net371;
wire net372_c1;
wire net372;
wire net373_c1;
wire net373;
wire net374_c1;
wire net374;
wire net375_c1;
wire net375;
wire net376_c1;
wire net376;
wire net377_c1;
wire net377;
wire net378_c1;
wire net378;
wire net379_c1;
wire net379;
wire net380_c1;
wire net380;
wire net381_c1;
wire net381;
wire net382_c1;
wire net382;
wire net383_c1;
wire net383;
wire net384_c1;
wire net384;
wire net385_c1;
wire net385;
wire net386_c1;
wire net386;
wire net387_c1;
wire net387;
wire net388_c1;
wire net388;
wire net389_c1;
wire net389;
wire net390_c1;
wire net390;
wire net391_c1;
wire net391;
wire net392_c1;
wire net392;
wire net393_c1;
wire net393;
wire net394_c1;
wire net394;
wire net395_c1;
wire net395;
wire net396_c1;
wire net396;
wire net397_c1;
wire net397;
wire net398_c1;
wire net398;
wire net399_c1;
wire net399;
wire net400_c1;
wire net400;
wire net401_c1;
wire net401;
wire net402_c1;
wire net402;
wire net403_c1;
wire net403;
wire net404_c1;
wire net404;
wire net405_c1;
wire net405;
wire net406_c1;
wire net406;
wire net407_c1;
wire net407;
wire net408_c1;
wire net408;
wire net409_c1;
wire net409;
wire net410_c1;
wire net410;
wire net411_c1;
wire net411;
wire net412_c1;
wire net412;
wire net413_c1;
wire net413;
wire net414_c1;
wire net414;
wire net415_c1;
wire net415;
wire net416_c1;
wire net416;
wire net417_c1;
wire net417;
wire net418_c1;
wire net418;
wire net419_c1;
wire net419;
wire net420_c1;
wire net420;
wire net421_c1;
wire net421;
wire net422_c1;
wire net422;
wire net423_c1;
wire net423;
wire net424_c1;
wire net424;
wire net425_c1;
wire net425;
wire net426_c1;
wire net426;
wire net427_c1;
wire net427;
wire net428_c1;
wire net428;
wire net429_c1;
wire net429;
wire net430_c1;
wire net430;
wire net431_c1;
wire net431;
wire net432_c1;
wire net432;
wire net433_c1;
wire net433;
wire net434_c1;
wire net434;
wire net435_c1;
wire net435;
wire net436_c1;
wire net436;
wire net437_c1;
wire net437;
wire net438_c1;
wire net438;
wire net439_c1;
wire net439;
wire net440_c1;
wire net440;
wire net441_c1;
wire net441;
wire net442_c1;
wire net442;
wire net443_c1;
wire net443;
wire net444_c1;
wire net444;
wire net445_c1;
wire net445;
wire net446_c1;
wire net446;
wire net447_c1;
wire net447;
wire net448_c1;
wire net448;
wire net449_c1;
wire net449;
wire net450_c1;
wire net450;
wire net451_c1;
wire net451;
wire net452_c1;
wire net452;
wire net453_c1;
wire net453;
wire net454_c1;
wire net454;
wire net455_c1;
wire net455;
wire net456_c1;
wire net456;
wire net457_c1;
wire net457;
wire net458_c1;
wire net458;
wire net459_c1;
wire net459;
wire net460_c1;
wire net460;
wire net461_c1;
wire net461;
wire net462_c1;
wire net462;
wire net463_c1;
wire net463;
wire net464_c1;
wire net464;
wire net465_c1;
wire net465;
wire net466_c1;
wire net466;
wire net467_c1;
wire net467;
wire net468_c1;
wire net468;
wire net469_c1;
wire net469;
wire net470_c1;
wire net470;
wire net471_c1;
wire net471;
wire net472_c1;
wire net472;
wire net473_c1;
wire net473;
wire net474_c1;
wire net474;
wire net475_c1;
wire net475;
wire net476_c1;
wire net476;
wire net477_c1;
wire net477;
wire net478_c1;
wire net478;
wire net479_c1;
wire net479;
wire net480_c1;
wire net480;
wire net481_c1;
wire net481;
wire net482_c1;
wire net482;
wire net483_c1;
wire net483;
wire net484_c1;
wire net484;
wire net485_c1;
wire net485;
wire net486_c1;
wire net486;
wire net487_c1;
wire net487;
wire net488_c1;
wire net488;
wire net489_c1;
wire net489;
wire net490_c1;
wire net490;
wire net491_c1;
wire net491;
wire net492_c1;
wire net492;
wire net493_c1;
wire net493;
wire net494_c1;
wire net494;
wire net495_c1;
wire net495;
wire net496_c1;
wire net496;
wire net497_c1;
wire net497;
wire net498_c1;
wire net498;
wire net499_c1;
wire net499;
wire net500_c1;
wire net500;
wire net501_c1;
wire net501;
wire net502_c1;
wire net502;
wire net503_c1;
wire net503;
wire net504_c1;
wire net504;
wire net505_c1;
wire net505;
wire net506_c1;
wire net506;
wire net507_c1;
wire net507;
wire net508_c1;
wire net508;
wire net509_c1;
wire net509;
wire net510_c1;
wire net510;
wire net511_c1;
wire net511;
wire net512_c1;
wire net512;
wire net513_c1;
wire net513;
wire net514_c1;
wire net514;
wire net515_c1;
wire net515;
wire net516_c1;
wire net516;
wire net517_c1;
wire net517;
wire net518_c1;
wire net518;
wire net519_c1;
wire net519;
wire net520_c1;
wire net520;
wire net521_c1;
wire net521;
wire net522_c1;
wire net522;
wire net523_c1;
wire net523;
wire net524_c1;
wire net524;
wire net525_c1;
wire net525;
wire net526_c1;
wire net526;
wire net527_c1;
wire net527;
wire net528_c1;
wire net528;
wire net529_c1;
wire net529;
wire net530_c1;
wire net530;
wire net531_c1;
wire net531;
wire net532_c1;
wire net532;
wire net533_c1;
wire net533;
wire net534_c1;
wire net534;
wire net535_c1;
wire net535;
wire net536_c1;
wire net536;
wire net537_c1;
wire net537;
wire net538_c1;
wire net538;
wire net539_c1;
wire net539;
wire net540_c1;
wire net540;
wire net541_c1;
wire net541;
wire net542_c1;
wire net542;
wire net543_c1;
wire net543;
wire net544_c1;
wire net544;
wire net545_c1;
wire net545;
wire net546_c1;
wire net546;
wire net547_c1;
wire net547;
wire net548_c1;
wire net548;
wire net549_c1;
wire net549;
wire net550_c1;
wire net550;
wire net551_c1;
wire net551;
wire net552_c1;
wire net552;
wire net553_c1;
wire net553;
wire net554_c1;
wire net554;
wire net555_c1;
wire net555;
wire net556_c1;
wire net556;
wire net557_c1;
wire net557;
wire net558_c1;
wire net558;
wire net559_c1;
wire net559;
wire net560_c1;
wire net560;
wire net561_c1;
wire net561;
wire net562_c1;
wire net562;
wire net563_c1;
wire net563;
wire net564_c1;
wire net564;
wire net565_c1;
wire net565;
wire net566_c1;
wire net566;
wire net567_c1;
wire net567;
wire net568_c1;
wire net568;
wire net569_c1;
wire net569;
wire net570_c1;
wire net570;
wire net571_c1;
wire net571;
wire net572_c1;
wire net572;
wire net573_c1;
wire net573;
wire net574_c1;
wire net574;
wire net575_c1;
wire net575;
wire net576_c1;
wire net576;
wire net577_c1;
wire net577;
wire net578_c1;
wire net578;
wire net579_c1;
wire net579;
wire net580_c1;
wire net580;
wire net581_c1;
wire net581;
wire net582_c1;
wire net582;
wire net583_c1;
wire net583;
wire net584_c1;
wire net584;
wire net585_c1;
wire net585;
wire net586_c1;
wire net586;
wire net587_c1;
wire net587;
wire net588_c1;
wire net588;
wire net589_c1;
wire net589;
wire net590_c1;
wire net590;
wire net591_c1;
wire net591;
wire net592_c1;
wire net592;
wire net593_c1;
wire net593;
wire net594_c1;
wire net594;
wire net595_c1;
wire net595;
wire net596_c1;
wire net596;
wire net597_c1;
wire net597;
wire net598_c1;
wire net598;
wire net599_c1;
wire net599;
wire net600_c1;
wire net600;
wire net601_c1;
wire net601;
wire net602_c1;
wire net602;
wire net603_c1;
wire net603;
wire net604_c1;
wire net604;
wire net605_c1;
wire net605;
wire net606_c1;
wire net606;
wire net607_c1;
wire net607;
wire net608_c1;
wire net608;
wire net609_c1;
wire net609;
wire net610_c1;
wire net610;
wire net611_c1;
wire net611;
wire net612_c1;
wire net612;
wire net613_c1;
wire net613;
wire net614_c1;
wire net614;
wire net615_c1;
wire net615;
wire net616_c1;
wire net616;
wire net617_c1;
wire net617;
wire net618_c1;
wire net618;
wire net619_c1;
wire net619;
wire net620_c1;
wire net620;
wire net621_c1;
wire net621;
wire net622_c1;
wire net622;
wire net623_c1;
wire net623;
wire net624_c1;
wire net624;
wire net625_c1;
wire net625;
wire net626_c1;
wire net626;
wire net627_c1;
wire net627;
wire net628_c1;
wire net628;
wire net629_c1;
wire net629;
wire net630_c1;
wire net630;
wire net631_c1;
wire net631;
wire net632_c1;
wire net632;
wire net633_c1;
wire net633;
wire net634_c1;
wire net634;
wire net635_c1;
wire net635;
wire net636_c1;
wire net636;
wire net637_c1;
wire net637;
wire net638_c1;
wire net638;
wire net639_c1;
wire net639;
wire net640_c1;
wire net640;
wire net641_c1;
wire net641;
wire net642_c1;
wire net642;
wire net643_c1;
wire net643;
wire net644_c1;
wire net644;
wire net645_c1;
wire net645;
wire net646_c1;
wire net646;
wire net647_c1;
wire net647;
wire net648_c1;
wire net648;
wire net649_c1;
wire net649;
wire net650_c1;
wire net650;
wire net651_c1;
wire net651;
wire net652_c1;
wire net652;
wire net653_c1;
wire net653;
wire net654_c1;
wire net654;
wire net655_c1;
wire net655;
wire net656_c1;
wire net656;
wire net657_c1;
wire net657;
wire net658_c1;
wire net658;
wire net659_c1;
wire net659;
wire net660_c1;
wire net660;
wire net661_c1;
wire net661;
wire net662_c1;
wire net662;
wire net663_c1;
wire net663;
wire net664_c1;
wire net664;
wire net665_c1;
wire net665;
wire net666_c1;
wire net666;
wire net667_c1;
wire net667;
wire net668_c1;
wire net668;
wire net669_c1;
wire net669;
wire net670_c1;
wire net670;
wire net671_c1;
wire net671;
wire net672_c1;
wire net672;
wire net673_c1;
wire net673;
wire net674_c1;
wire net674;
wire net675_c1;
wire net675;
wire net676_c1;
wire net676;
wire net677_c1;
wire net677;
wire net678_c1;
wire net678;
wire net679_c1;
wire net679;
wire net680_c1;
wire net680;
wire net681_c1;
wire net681;
wire net682_c1;
wire net682;
wire net683_c1;
wire net683;
wire net684_c1;
wire net684;
wire net685_c1;
wire net685;
wire net686_c1;
wire net686;
wire net687_c1;
wire net687;
wire net688_c1;
wire net688;
wire net689_c1;
wire net689;
wire net690_c1;
wire net690;
wire net691_c1;
wire net691;
wire net692_c1;
wire net692;
wire net693_c1;
wire net693;
wire net694_c1;
wire net694;
wire net695_c1;
wire net695;
wire net696_c1;
wire net696;
wire net697_c1;
wire net697;
wire net698_c1;
wire net698;
wire net699_c1;
wire net699;
wire net700_c1;
wire net700;
wire net701_c1;
wire net701;
wire net702_c1;
wire net702;
wire net703_c1;
wire net703;
wire net704_c1;
wire net704;
wire net705_c1;
wire net705;
wire net706_c1;
wire net706;
wire net707_c1;
wire net707;
wire net708_c1;
wire net708;
wire net709_c1;
wire net709;
wire net710_c1;
wire net710;
wire net711_c1;
wire net711;
wire net712_c1;
wire net712;
wire net713_c1;
wire net713;
wire net714_c1;
wire net714;
wire net715_c1;
wire net715;
wire net716_c1;
wire net716;
wire net717_c1;
wire net717;
wire net718_c1;
wire net718;
wire net719_c1;
wire net719;
wire net720_c1;
wire net720;
wire net721_c1;
wire net721;
wire net722_c1;
wire net722;
wire net723_c1;
wire net723;
wire net724_c1;
wire net724;
wire net725_c1;
wire net725;
wire net726_c1;
wire net726;
wire net727_c1;
wire net727;
wire net728_c1;
wire net728;
wire net729_c1;
wire net729;
wire net730_c1;
wire net730;
wire net731_c1;
wire net731;
wire net732_c1;
wire net732;
wire net733_c1;
wire net733;
wire net734_c1;
wire net734;
wire net735_c1;
wire net735;
wire net736_c1;
wire net736;
wire net737_c1;
wire net737;
wire net738_c1;
wire net738;
wire net739_c1;
wire net739;
wire net740_c1;
wire net740;
wire net741_c1;
wire net741;
wire net742_c1;
wire net742;
wire net743_c1;
wire net743;
wire net744_c1;
wire net744;
wire net745_c1;
wire net745;
wire net746_c1;
wire net746;
wire net747_c1;
wire net747;
wire net748_c1;
wire net748;
wire net749_c1;
wire net749;
wire net750_c1;
wire net750;
wire net751_c1;
wire net751;
wire net752_c1;
wire net752;
wire net753_c1;
wire net753;
wire net754_c1;
wire net754;
wire net755_c1;
wire net755;
wire net756_c1;
wire net756;
wire net757_c1;
wire net757;
wire net758_c1;
wire net758;
wire net759_c1;
wire net759;
wire net760_c1;
wire net760;
wire net761_c1;
wire net761;
wire net762_c1;
wire net762;
wire net763_c1;
wire net763;
wire net764_c1;
wire net764;
wire net765_c1;
wire net765;
wire net766_c1;
wire net766;
wire net767_c1;
wire net767;
wire net768_c1;
wire net768;
wire net769_c1;
wire net769;
wire net770_c1;
wire net770;
wire net771_c1;
wire net771;
wire net772_c1;
wire net772;
wire net773_c1;
wire net773;
wire net774_c1;
wire net774;
wire net775_c1;
wire net775;
wire net776_c1;
wire net776;
wire net777_c1;
wire net777;
wire net778_c1;
wire net778;
wire net779_c1;
wire net779;
wire net780_c1;
wire net780;
wire net781_c1;
wire net781;
wire net782_c1;
wire net782;
wire net783_c1;
wire net783;
wire net784_c1;
wire net784;
wire net785_c1;
wire net785;
wire net786_c1;
wire net786;
wire net787_c1;
wire net787;
wire net788_c1;
wire net788;
wire net789_c1;
wire net789;
wire net790_c1;
wire net790;
wire net791_c1;
wire net791;
wire net792_c1;
wire net792;
wire net793_c1;
wire net793;
wire net794_c1;
wire net794;
wire net795_c1;
wire net795;
wire net796_c1;
wire net796;
wire net797_c1;
wire net797;
wire net798_c1;
wire net798;
wire net799_c1;
wire net799;
wire net800_c1;
wire net800;
wire net801_c1;
wire net801;
wire net802_c1;
wire net802;
wire net803_c1;
wire net803;
wire net804_c1;
wire net804;
wire net805_c1;
wire net805;
wire net806_c1;
wire net806;
wire net807_c1;
wire net807;
wire net808_c1;
wire net808;
wire net809_c1;
wire net809;
wire net810_c1;
wire net810;
wire net811_c1;
wire net811;
wire net812_c1;
wire net812;
wire net813_c1;
wire net813;
wire net814_c1;
wire net814;
wire net815_c1;
wire net815;
wire net816_c1;
wire net816;
wire net817_c1;
wire net817;
wire net818_c1;
wire net818;
wire net819_c1;
wire net819;
wire net820_c1;
wire net820;
wire net821_c1;
wire net821;
wire net822_c1;
wire net822;
wire net823_c1;
wire net823;
wire net824_c1;
wire net824;
wire net825_c1;
wire net825;
wire net826_c1;
wire net826;
wire net827_c1;
wire net827;
wire net828_c1;
wire net828;
wire net829_c1;
wire net829;
wire net830_c1;
wire net830;
wire net831_c1;
wire net831;
wire net832_c1;
wire net832;
wire net833_c1;
wire net833;
wire net834_c1;
wire net834;
wire net835_c1;
wire net835;
wire net836_c1;
wire net836;
wire net837_c1;
wire net837;
wire net838_c1;
wire net838;
wire net839_c1;
wire net839;
wire net840_c1;
wire net840;
wire net841_c1;
wire net841;
wire net842_c1;
wire net842;
wire net843_c1;
wire net843;
wire net844_c1;
wire net844;
wire net845_c1;
wire net845;
wire net846_c1;
wire net846;
wire net847_c1;
wire net847;
wire net848_c1;
wire net848;
wire net849_c1;
wire net849;
wire net850_c1;
wire net850;
wire net851_c1;
wire net851;
wire net852_c1;
wire net852;
wire net853_c1;
wire net853;
wire net854_c1;
wire net854;
wire net855_c1;
wire net855;
wire net856_c1;
wire net856;
wire net857_c1;
wire net857;
wire net858_c1;
wire net858;
wire net859_c1;
wire net859;
wire net860_c1;
wire net860;
wire net861_c1;
wire net861;
wire net862_c1;
wire net862;
wire net863_c1;
wire net863;
wire net864_c1;
wire net864;
wire net865_c1;
wire net865;
wire net866_c1;
wire net866;
wire net867_c1;
wire net867;
wire net868_c1;
wire net868;
wire net869_c1;
wire net869;
wire net870_c1;
wire net870;
wire net871_c1;
wire net871;
wire net872_c1;
wire net872;
wire net873_c1;
wire net873;
wire net874_c1;
wire net874;
wire net875_c1;
wire net875;
wire net876_c1;
wire net876;
wire net877_c1;
wire net877;
wire net878_c1;
wire net878;
wire net879_c1;
wire net879;
wire net880_c1;
wire net880;
wire net881_c1;
wire net881;
wire net882_c1;
wire net882;
wire net883_c1;
wire net883;
wire net884_c1;
wire net884;
wire net885_c1;
wire net885;
wire net886_c1;
wire net886;
wire net887_c1;
wire net887;
wire net888_c1;
wire net888;
wire net889_c1;
wire net889;
wire net890_c1;
wire net890;
wire net891_c1;
wire net891;
wire net892_c1;
wire net892;
wire net893_c1;
wire net893;
wire net894_c1;
wire net894;
wire net895_c1;
wire net895;
wire net896_c1;
wire net896;
wire net897_c1;
wire net897;
wire net898_c1;
wire net898;
wire net899_c1;
wire net899;
wire net900_c1;
wire net900;
wire net901_c1;
wire net901;
wire net902_c1;
wire net902;
wire net903_c1;
wire net903;
wire net904_c1;
wire net904;
wire net905_c1;
wire net905;
wire net906_c1;
wire net906;
wire net907_c1;
wire net907;
wire net908_c1;
wire net908;
wire net909_c1;
wire net909;
wire net910_c1;
wire net910;
wire net911_c1;
wire net911;
wire net912_c1;
wire net912;
wire net913_c1;
wire net913;
wire net914_c1;
wire net914;
wire net915_c1;
wire net915;
wire net916_c1;
wire net916;
wire net917_c1;
wire net917;
wire net918_c1;
wire net918;
wire net919_c1;
wire net919;
wire net920_c1;
wire net920;
wire net921_c1;
wire net921;
wire net922_c1;
wire net922;
wire net923_c1;
wire net923;
wire net924_c1;
wire net924;
wire net925_c1;
wire net925;
wire net926_c1;
wire net926;
wire net927_c1;
wire net927;
wire net928_c1;
wire net928;
wire net929_c1;
wire net929;
wire net930_c1;
wire net930;
wire net931_c1;
wire net931;
wire net932_c1;
wire net932;
wire net933_c1;
wire net933;
wire net934_c1;
wire net934;
wire net935_c1;
wire net935;
wire net936_c1;
wire net936;
wire net937_c1;
wire net937;
wire net938_c1;
wire net938;
wire net939_c1;
wire net939;
wire net940_c1;
wire net940;
wire net941_c1;
wire net941;
wire net942_c1;
wire net942;
wire net943_c1;
wire net943;
wire net944_c1;
wire net944;
wire net945_c1;
wire net945;
wire net946_c1;
wire net946;
wire net947_c1;
wire net947;
wire net948_c1;
wire net948;
wire net949_c1;
wire net949;
wire net950_c1;
wire net950;
wire net951_c1;
wire net951;
wire net952_c1;
wire net952;
wire net953_c1;
wire net953;
wire net954_c1;
wire net954;
wire net955_c1;
wire net955;
wire net956_c1;
wire net956;
wire net957_c1;
wire net957;
wire net958_c1;
wire net958;
wire net959_c1;
wire net959;
wire net960_c1;
wire net960;
wire net961_c1;
wire net961;
wire net962_c1;
wire net962;
wire net963_c1;
wire net963;
wire net964_c1;
wire net964;
wire net965_c1;
wire net965;
wire net966_c1;
wire net966;
wire net967_c1;
wire net967;
wire net968_c1;
wire net968;
wire net969_c1;
wire net969;
wire net970_c1;
wire net970;
wire net971_c1;
wire net971;
wire net972_c1;
wire net972;
wire net973_c1;
wire net973;
wire net974_c1;
wire net974;
wire net975_c1;
wire net975;
wire net976_c1;
wire net976;
wire net977_c1;
wire net977;
wire net978_c1;
wire net978;
wire net979_c1;
wire net979;
wire net980_c1;
wire net980;
wire net981_c1;
wire net981;
wire net982_c1;
wire net982;
wire net983_c1;
wire net983;
wire net984_c1;
wire net984;
wire net985_c1;
wire net985;
wire net986_c1;
wire net986;
wire net987_c1;
wire net987;
wire net988_c1;
wire net988;
wire net989_c1;
wire net989;
wire net990_c1;
wire net990;
wire net991_c1;
wire net991;
wire net992_c1;
wire net992;
wire net993_c1;
wire net993;
wire net994_c1;
wire net994;
wire net995_c1;
wire net995;
wire net996_c1;
wire net996;
wire net997_c1;
wire net997;
wire net998_c1;
wire net998;
wire net999_c1;
wire net999;
wire net1000_c1;
wire net1000;
wire net1001_c1;
wire net1001;
wire net1002_c1;
wire net1002;
wire net1003_c1;
wire net1003;
wire net1004_c1;
wire net1004;
wire net1005_c1;
wire net1005;
wire net1006_c1;
wire net1006;
wire GCLK_Pad;
wire net1007;
wire net1008_c1;
wire net1008;

DFFT DFFT_199__FPB_n526(net967,net362,net440_c1);
XOR2T XOR2T_29_n41(net777,net355,net484,net12_c1);
AND2T AND2T_110_n122(net985,net210,net478,net99_c1);
AND2T AND2T_102_n114(net851,net300,net455,net100_c1);
AND2T AND2T_103_n115(net837,net100,net278,net104_c1);
AND2T AND2T_120_n132(net845,net173,net487,net107_c1);
AND2T AND2T_112_n124(net751,net180,net488,net108_c1);
AND2T AND2T_104_n116(net813,net289,net461,net109_c1);
AND2T AND2T_121_n133(net849,net107,net154,net112_c1);
AND2T AND2T_113_n125(net565,net29,net450,net113_c1);
AND2T AND2T_122_n134(net835,net161,net492,net117_c1);
AND2T AND2T_114_n126(net687,net337,net454,net118_c1);
AND2T AND2T_106_n118(net937,net372,net473,net119_c1);
AND2T AND2T_123_n135(net1003,net166,net465,net121_c1);
AND2T AND2T_107_n119(net959,net119,net33,net123_c1);
AND2T AND2T_124_n136(net989,net209,net477,net125_c1);
AND2T AND2T_133_n145(net873,net124,net120,net128_c1);
AND2T AND2T_125_n137(net905,net132,net483,net129_c1);
AND2T AND2T_134_n161(net633,net10,net30,net127_c1);
AND2T AND2T_119_n131(net601,net98,net114,net102_c1);
AND2T AND2T_135_n162(net587,net238,net501,net131_c1);
AND2T AND2T_136_n163(net510,net15,net472,net133_c1);
AND2T AND2T_137_n164(net771,net399,net260,net135_c1);
AND2T AND2T_4_n16(net567,net284,net391,net11_c1);
AND2T AND2T_7_n19(net543,net352,net348,net25_c1);
AND2T AND2T_8_n20(net509,net374,net485,net2_c1);
OR2T OR2T_9_n21(net535,net251,net176,net3_c1);
NOTT NOTT_5_n17(net523,net298,net15_c1);
NOTT NOTT_6_n18(net583,net373,net20_c1);
AND2T AND2T_22_n34(net603,net13,net6,net18_c1);
AND2T AND2T_31_n43(net625,net28,net493,net22_c1);
AND2T AND2T_23_n35(net602,net18,net24,net23_c1);
AND2T AND2T_15_n27(net597,net19,net498,net24_c1);
AND2T AND2T_40_n52(net568,net21,net50,net27_c1);
AND2T AND2T_24_n36(net529,net363,net475,net29_c1);
AND2T AND2T_41_n53(net611,net27,net44,net32_c1);
AND2T AND2T_33_n45(net789,net229,net497,net33_c1);
AND2T AND2T_25_n37(net659,net358,net211,net34_c1);
AND2T AND2T_17_n29(net631,net367,net384,net35_c1);
AND2T AND2T_50_n62(net632,net245,net418,net37_c1);
AND2T AND2T_34_n46(net634,net322,net340,net39_c1);
AND2T AND2T_51_n63(net657,net283,net250,net42_c1);
AND2T AND2T_27_n39(net899,net343,net480,net45_c1);
AND2T AND2T_28_n40(net719,net268,net12,net8_c1);
AND2T AND2T_60_n72(net665,net41,net64,net47_c1);
AND2T AND2T_61_n73(net713,net142,net230,net52_c1);
AND2T AND2T_45_n57(net588,net49,net43,net54_c1);
AND2T AND2T_37_n49(net778,net386,net387,net55_c1);
AND2T AND2T_38_n50(net551,net341,net338,net16_c1);
AND2T AND2T_62_n74(net688,net318,net413,net58_c1);
AND2T AND2T_54_n66(net997,net292,net410,net59_c1);
AND2T AND2T_46_n58(net791,net274,net65,net60_c1);
AND2T AND2T_63_n75(net573,net35,net417,net63_c1);
AND2T AND2T_47_n59(net815,net291,net411,net65_c1);
AND2T AND2T_48_n60(net814,net281,net414,net26_c1);
AND2T AND2T_72_n84(net508,net329,net447,net67_c1);
AND2T AND2T_64_n76(net900,net365,net421,net68_c1);
AND2T AND2T_56_n68(net645,net216,net326,net69_c1);
AND2T AND2T_65_n77(net921,net68,net198,net72_c1);
AND2T AND2T_57_n69(net571,net156,net426,net73_c1);
AND2T AND2T_74_n86(net646,net364,net452,net75_c1);
AND2T AND2T_83_n95(net819,net74,net62,net77_c1);
AND2T AND2T_75_n87(net707,net287,net204,net78_c1);
AND2T AND2T_84_n96(net721,net269,net205,net80_c1);
AND2T AND2T_85_n97(net705,net162,net236,net82_c1);
AND2T AND2T_87_n99(net943,net296,net435,net85_c1);
OR2T OR2T_10_n22(net574,net159,net265,net5_c1);
OR2T OR2T_11_n23(net530,net353,net339,net7_c1);
OR2T OR2T_20_n32(net617,net259,net469,net9_c1);
OR2T OR2T_21_n33(net589,net375,net239,net13_c1);
OR2T OR2T_13_n25(net541,net232,net490,net14_c1);
OR2T OR2T_30_n42(net714,net383,net489,net17_c1);
OR2T OR2T_14_n26(net590,net359,net494,net19_c1);
OR2T OR2T_18_n30(net775,net225,net463,net4_c1);
OR2T OR2T_26_n38(net660,net34,net0,net40_c1);
OR2T OR2T_19_n31(net776,net4,net333,net6_c1);
OR2T OR2T_43_n55(net544,net282,net366,net43_c1);
OR2T OR2T_52_n64(net559,net42,net423,net48_c1);
OR2T OR2T_44_n56(net553,net158,net502,net49_c1);
OR2T OR2T_36_n48(net612,net249,net500,net50_c1);
OR2T OR2T_53_n65(net706,net48,net427,net53_c1);
OR2T OR2T_70_n82(net961,net51,net436,net57_c1);
OR2T OR2T_71_n83(net821,net57,net305,net62_c1);
OR2T OR2T_55_n67(net711,net258,net422,net64_c1);
OR2T OR2T_80_n92(net973,net168,net457,net66_c1);
OR2T OR2T_81_n93(net953,net314,net301,net70_c1);
OR2T OR2T_73_n85(net658,net290,net297,net71_c1);
OR2T OR2T_58_n70(net673,net303,net437,net36_c1);
OR2T OR2T_82_n94(net859,net181,net420,net74_c1);
OR2T OR2T_66_n78(net651,net285,net323,net76_c1);
OR2T OR2T_59_n71(net663,net36,net442,net41_c1);
OR2T OR2T_67_n79(net664,net76,net425,net79_c1);
OR2T OR2T_68_n80(net675,net79,net432,net46_c1);
OR2T OR2T_76_n88(net649,net295,net75,net81_c1);
OR2T OR2T_69_n81(net735,net46,net47,net51_c1);
OR2T OR2T_77_n89(net652,net81,net71,net83_c1);
OR2T OR2T_78_n90(net708,net149,net83,net56_c1);
OR2T OR2T_86_n98(net913,net336,net80,net84_c1);
OR2T OR2T_79_n91(net650,net197,net182,net61_c1);
NOTT NOTT_12_n24(net627,net288,net10_c1);
NOTT NOTT_32_n44(net720,net273,net28_c1);
NOTT NOTT_16_n28(net805,net276,net30_c1);
NOTT NOTT_42_n54(net527,net215,net38_c1);
NOTT NOTT_35_n47(net613,net294,net44_c1);
NOTT NOTT_39_n51(net554,net270,net21_c1);
NOTT NOTT_49_n61(net681,net356,net31_c1);
OR2T OR2T_100_n112(net954,net90,net110,net93_c1);
OR2T OR2T_101_n113(net955,net93,net479,net96_c1);
OR2T OR2T_111_n123(net975,net99,net306,net103_c1);
OR2T OR2T_105_n117(net799,net327,net467,net114_c1);
OR2T OR2T_130_n142(net999,net111,net491,net116_c1);
OR2T OR2T_131_n143(net879,net312,net496,net120_c1);
OR2T OR2T_115_n127(net749,net118,net108,net122_c1);
OR2T OR2T_108_n120(net725,net123,net192,net92_c1);
OR2T OR2T_132_n144(net867,net187,net499,net124_c1);
OR2T OR2T_116_n128(net935,net122,net103,net126_c1);
OR2T OR2T_109_n121(net727,net92,net380,net95_c1);
OR2T OR2T_117_n129(net923,net126,net460,net130_c1);
OR2T OR2T_118_n130(net604,net202,net466,net98_c1);
OR2T OR2T_126_n138(net907,net377,net217,net132_c1);
OR2T OR2T_127_n139(net897,net129,net163,net134_c1);
OR2T OR2T_128_n140(net927,net134,net302,net106_c1);
OR2T OR2T_129_n141(net998,net106,net486,net111_c1);
OR2T OR2T_139_n166(net914,net310,net174,net139_c1);
AND2T AND2T_94_n106(net968,net97,net330,net101_c1);
AND2T AND2T_95_n107(net976,net191,net445,net105_c1);
AND2T AND2T_88_n100(net736,net167,net441,net86_c1);
AND2T AND2T_96_n108(net956,net105,net203,net110_c1);
AND2T AND2T_89_n101(net898,net143,net446,net87_c1);
AND2T AND2T_97_n109(net852,net169,net468,net115_c1);
AND2T AND2T_98_n110(net874,net115,net148,net88_c1);
AND2T AND2T_99_n111(net861,net157,net474,net90_c1);
DFFT DFFT_200__FPB_n527(net969,net440,net447_c1);
DFFT DFFT_201__FPB_n528(net618,net346,net452_c1);
DFFT DFFT_210__FPB_n537(net737,net172,net456_c1);
DFFT DFFT_202__FPB_n529(net974,net179,net457_c1);
DFFT DFFT_203__FPB_n530(net862,net335,net420_c1);
DFFT DFFT_211__FPB_n538(net983,net85,net462_c1);
DFFT DFFT_204__FPB_n531(net695,net243,net424_c1);
DFFT DFFT_220__FPB_n547(net875,net459,net468_c1);
DFFT DFFT_212__FPB_n539(net696,net235,net464_c1);
DFFT DFFT_213__FPB_n540(net741,net464,net428_c1);
DFFT DFFT_205__FPB_n532(net757,net424,net429_c1);
DFFT DFFT_221__FPB_n548(net850,net88,net474_c1);
DFFT DFFT_150__FBL_n477(net908,net190,net403_c1);
DFFT DFFT_214__FPB_n541(net743,net428,net433_c1);
DFFT DFFT_206__FPB_n533(net941,net429,net435_c1);
DFFT DFFT_230__FPB_n557(net960,net147,net478_c1);
DFFT DFFT_222__FPB_n549(net970,net101,net479_c1);
DFFT DFFT_151__FBL_n478(net880,net320,net404_c1);
DFFT DFFT_143__FPB_n185(net679,net201,net416_c1);
DFFT DFFT_223__FPB_n550(net783,net385,net438_c1);
DFFT DFFT_215__FPB_n542(net744,net433,net439_c1);
DFFT DFFT_207__FPB_n534(net689,net275,net441_c1);
DFFT DFFT_231__FPB_n558(net929,net248,net482_c1);
DFFT DFFT_152__FBL_n479(net507,net224,net405_c1);
OR2T OR2T_90_n102(net924,net155,net307,net89_c1);
OR2T OR2T_91_n103(net922,net89,net451,net91_c1);
OR2T OR2T_92_n104(net738,net91,net456,net94_c1);
OR2T OR2T_93_n105(net984,net94,net462,net97_c1);
DFFT DFFT_144__FPB_n186(net742,net319,net419_c1);
DFFT DFFT_224__FPB_n551(net785,net438,net443_c1);
DFFT DFFT_216__FPB_n543(net986,net439,net445_c1);
DFFT DFFT_208__FPB_n535(net722,net299,net446_c1);
DFFT DFFT_240__FPB_n567(net846,net481,net487_c1);
DFFT DFFT_232__FPB_n559(net928,net482,net488_c1);
DFFT DFFT_160__FPB_n487(net536,net304,net490_c1);
DFFT DFFT_153__FBL_n480(net595,net195,net392_c1);
DFFT DFFT_145__FBL_n472(net822,net331,net393_c1);
DFFT DFFT_233__FPB_n560(net552,net332,net450_c1);
DFFT DFFT_225__FPB_n552(net786,net443,net448_c1);
DFFT DFFT_217__FPB_n544(net881,net234,net449_c1);
DFFT DFFT_209__FPB_n536(net728,net313,net451_c1);
DFFT DFFT_241__FPB_n568(net836,net112,net492_c1);
DFFT DFFT_161__FPB_n488(net614,net247,net494_c1);
DFFT DFFT_154__FBL_n481(net537,net308,net395_c1);
DFFT DFFT_146__FBL_n473(net911,net315,net394_c1);
DFFT DFFT_234__FPB_n561(net682,net309,net454_c1);
DFFT DFFT_226__FPB_n553(net843,net448,net455_c1);
DFFT DFFT_218__FPB_n545(net882,net449,net453_c1);
DFFT DFFT_250__FPB_n577(net1005,net116,net496_c1);
DFFT DFFT_242__FPB_n569(net755,net378,net495_c1);
DFFT DFFT_170__FPB_n497(net792,net261,net497_c1);
DFFT DFFT_162__FPB_n489(net542,net1008,net498_c1);
DFFT DFFT_155__FBL_n482(net784,net316,net396_c1);
DFFT DFFT_147__FBL_n474(net584,net350,net397_c1);
DFFT DFFT_243__FPB_n570(net756,net495,net458_c1);
DFFT DFFT_235__FPB_n562(net936,net95,net460_c1);
DFFT DFFT_227__FPB_n554(net790,net104,net461_c1);
DFFT DFFT_219__FPB_n546(net876,net453,net459_c1);
DFFT DFFT_163__FPB_n490(net838,net379,net463_c1);
DFFT DFFT_251__FPB_n578(net868,net70,net499_c1);
DFFT DFFT_171__FPB_n498(net528,net218,net500_c1);
DFFT DFFT_156__FBL_n483(net807,net324,net398_c1);
DFFT DFFT_148__FBL_n475(net598,net321,net399_c1);
DFFT DFFT_180__FPB_n507(net619,net170,net427_c1);
DFFT DFFT_244__FPB_n571(net1004,net458,net465_c1);
DFFT DFFT_236__FPB_n563(net893,net130,net466_c1);
DFFT DFFT_228__FPB_n555(net801,net208,net467_c1);
DFFT DFFT_164__FPB_n491(net620,net164,net469_c1);
DFFT DFFT_252__FPB_n579(net596,net405,net501_c1);
DFFT DFFT_172__FPB_n499(net566,net231,net502_c1);
DFFT DFFT_157__FBL_n484(net865,net194,net400_c1);
DFFT DFFT_149__FBL_n476(net820,net200,net401_c1);
DFFT DFFT_173__FPB_n500(net628,net150,net406_c1);
DFFT DFFT_181__FPB_n508(net930,net237,net431_c1);
DFFT DFFT_253__FPB_n580(net772,net263,net472_c1);
DFFT DFFT_245__FPB_n572(net990,net253,net470_c1);
DFFT DFFT_237__FPB_n564(net831,net389,net471_c1);
DFFT DFFT_229__FPB_n556(net962,net394,net473_c1);
DFFT DFFT_165__FPB_n492(net524,net177,net475_c1);
DFFT DFFT_158__FBL_n485(net506,net178,net402_c1);
DFFT DFFT_174__FPB_n501(net800,net406,net407_c1);
DFFT DFFT_190__FPB_n517(net674,net430,net437_c1);
DFFT DFFT_182__FPB_n509(net942,net431,net434_c1);
DFFT DFFT_246__FPB_n573(net991,net470,net477_c1);
DFFT DFFT_238__FPB_n565(net832,net471,net476_c1);
DFFT DFFT_166__FPB_n493(net906,net357,net480_c1);
SPLITT Split_300_n627(net52,net185_c1,net313_c1);
SPLITT Split_301_n628(net185,net192_c1,net318_c1);
SPLITT Split_302_n629(net63,net197_c1,net323_c1);
SPLITT Split_310_n637(net77,net193_c1,net324_c1);
SPLITT Split_303_n630(net72,net155_c1,net285_c1);
SPLITT Split_311_n638(net193,net200_c1,net331_c1);
SPLITT Split_304_n631(net67,net163_c1,net290_c1);
SPLITT Split_312_n639(net82,net210_c1,net336_c1);
SPLITT Split_320_n647(net113,net209_c1,net337_c1);
SPLITT Split_305_n632(net78,net167_c1,net295_c1);
SPLITT Split_313_n640(net84,net166_c1,net296_c1);
SPLITT Split_321_n648(net102,net213_c1,net344_c1);
SPLITT Split_306_n633(net56,net174_c1,net301_c1);
SPLITT Split_314_n641(net86,net172_c1,net302_c1);
SPLITT Split_322_n649(net344,net224_c1,net350_c1);
SPLITT Split_330_n657(net131,net220_c1,net351_c1);
SPLITT Split_307_n634(net61,net179_c1,net306_c1);
SPLITT Split_315_n642(net87,net180_c1,net307_c1);
SPLITT Split_323_n650(net213,net178_c1,net308_c1);
SPLITT Split_331_n658(net351,net230_c1,net358_c1);
SPLITT Split_308_n635(net66,net186_c1,net310_c1);
SPLITT Split_316_n643(net96,net183_c1,net311_c1);
SPLITT Split_324_n651(net117,net187_c1,net312_c1);
SPLITT Split_260_n587(net221,net238_c1,net363_c1);
SPLITT Split_332_n659(net220,net236_c1,net364_c1);
SPLITT Split_340_n667(net354,net237_c1,net365_c1);
SPLITT Split_309_n636(net186,net191_c1,net314_c1);
SPLITT Split_317_n644(net311,net190_c1,net315_c1);
SPLITT Split_325_n652(net128,net189_c1,net316_c1);
SPLITT Split_333_n660(net133,net188_c1,net317_c1);
SPLITT Split_261_n588(net25,net242_c1,net370_c1);
SPLITT Split_341_n668(net226,net243_c1,net371_c1);
SPLITT Split_254_n581(net1,net196_c1,net319_c1);
SPLITT Split_318_n645(net183,net194_c1,net320_c1);
SPLITT Split_326_n653(net189,net195_c1,net321_c1);
SPLITT Split_334_n661(net317,net198_c1,net322_c1);
SPLITT Split_262_n589(net370,net250_c1,net374_c1);
SPLITT Split_270_n597(net244,net249_c1,net375_c1);
SPLITT Split_342_n669(net139,net246_c1,net376_c1);
SPLITT Split_350_n677(net233,net247_c1,net377_c1);
SPLITT Split_255_n582(net196,net201_c1,net325_c1);
SPLITT Split_263_n590(net242,net205_c1,net326_c1);
SPLITT Split_319_n646(net109,net202_c1,net327_c1);
SPLITT Split_327_n654(net127,net199_c1,net328_c1);
SPLITT Split_335_n662(net188,net204_c1,net329_c1);
SPLITT Split_343_n670(net376,net203_c1,net330_c1);
SPLITT Split_271_n598(net40,net255_c1,net380_c1);
SPLITT Split_351_n678(net140,net252_c1,net381_c1);
SPLITT Split_280_n607(net153,net161_c1,net289_c1);
SPLITT Split_256_n583(net11,net207_c1,net332_c1);
SPLITT Split_328_n655(net328,net211_c1,net333_c1);
SPLITT Split_336_n663(net135,net206_c1,net334_c1);
SPLITT Split_344_n671(net246,net208_c1,net335_c1);
SPLITT Split_272_n599(net255,net258_c1,net383_c1);
SPLITT Split_352_n679(net381,net259_c1,net384_c1);
SPLITT Split_360_n687(net397,net257_c1,net385_c1);
SPLITT Split_273_n600(net45,net141_c1,net267_c1);
SPLITT Split_281_n608(net39,net170_c1,net294_c1);
SPLITT Split_257_n584(net207,net214_c1,net338_c1);
SPLITT Split_265_n592(net3,net218_c1,net339_c1);
SPLITT Split_329_n656(net199,net216_c1,net340_c1);
SPLITT Split_337_n664(net334,net215_c1,net341_c1);
SPLITT Split_345_n672(net136,net212_c1,net342_c1);
SPLITT Split_353_n680(net252,net217_c1,net343_c1);
SPLITT Split_361_n688(net257,net260_c1,net387_c1);
DFFT DFFT_183__FPB_n510(net938,net434,net408_c1);
DFFT DFFT_175__FPB_n502(net806,net407,net409_c1);
SPLITT Split_274_n601(net267,net142_c1,net268_c1);
DFFT DFFT_191__FPB_n518(net712,net175,net442_c1);
SPLITT Split_282_n609(net55,net171_c1,net299_c1);
SPLITT Split_290_n617(net160,net173_c1,net300_c1);
DFFT DFFT_247__FPB_n574(net894,net171,net483_c1);
DFFT DFFT_239__FPB_n566(net844,net476,net481_c1);
DFFT DFFT_167__FPB_n494(net505,net254,net484_c1);
DFFT DFFT_159__FPB_n486(net557,net214,net485_c1);
SPLITT Split_258_n585(net20,net221_c1,net345_c1);
SPLITT Split_266_n593(net5,net222_c1,net346_c1);
SPLITT Split_338_n665(net206,net223_c1,net347_c1);
SPLITT Split_346_n673(net342,net225_c1,net348_c1);
SPLITT Split_354_n681(net416,net219_c1,net349_c1);
SPLITT Split_362_n689(net404,net262_c1,net388_c1);
SPLITT Split_370_n697(net256,net263_c1,net389_c1);
SPLITT Split_275_n602(net141,net143_c1,net269_c1);
SPLITT Split_283_n610(net16,net144_c1,net270_c1);
SPLITT Split_291_n618(net26,net181_c1,net305_c1);
SPLITT Split_259_n586(net345,net232_c1,net352_c1);
SPLITT Split_267_n594(net222,net231_c1,net353_c1);
SPLITT Split_339_n666(net137,net226_c1,net354_c1);
SPLITT Split_347_n674(net212,net229_c1,net355_c1);
SPLITT Split_355_n682(net349,net228_c1,net356_c1);
SPLITT Split_363_n690(net388,net227_c1,net357_c1);
SPLITT Split_371_n698(net398,net264_c1,net390_c1);
SPLITT Split_276_n603(net8,net146_c1,net271_c1);
SPLITT Split_284_n611(net32,net145_c1,net272_c1);
SPLITT Split_292_n619(net31,net184_c1,net309_c1);
SPLITT Split_268_n595(net14,net239_c1,net359_c1);
SPLITT Split_348_n675(net138,net233_c1,net360_c1);
SPLITT Split_356_n683(net219,net235_c1,net361_c1);
SPLITT Split_364_n691(net262,net234_c1,net362_c1);
SPLITT Split_372_n699(net390,net265_c1,net391_c1);
SPLITT Split_277_n604(net17,net149_c1,net273_c1);
SPLITT Split_285_n612(net272,net148_c1,net274_c1);
SPLITT Split_293_n620(net184,net147_c1,net275_c1);
SPLITT Split_373_n700(net264,net150_c1,net276_c1);
SPLITT Split_269_n596(net9,net244_c1,net366_c1);
SPLITT Split_349_n676(net360,net245_c1,net367_c1);
SPLITT Split_357_n684(net419,net241_c1,net368_c1);
SPLITT Split_365_n692(net392,net240_c1,net369_c1);
SPLITT Split_278_n605(net22,net153_c1,net277_c1);
SPLITT Split_286_n613(net145,net154_c1,net278_c1);
SPLITT Split_294_n621(net37,net152_c1,net279_c1);
SPLITT Split_374_n701(net400,net151_c1,net280_c1);
SPLITT Split_358_n685(net368,net248_c1,net372_c1);
SPLITT Split_366_n693(net369,net251_c1,net373_c1);
SPLITT Split_279_n606(net277,net157_c1,net281_c1);
SPLITT Split_287_n614(net38,net158_c1,net282_c1);
SPLITT Split_295_n622(net279,net156_c1,net283_c1);
SPLITT Split_375_n702(net280,net159_c1,net284_c1);
SPLITT Split_359_n686(net241,net253_c1,net378_c1);
SPLITT Split_367_n694(net240,net254_c1,net379_c1);
SPLITT Split_288_n615(net54,net160_c1,net286_c1);
SPLITT Split_296_n623(net152,net162_c1,net287_c1);
SPLITT Split_376_n703(net151,net164_c1,net288_c1);
SPLITT Split_368_n695(net396,net256_c1,net382_c1);
SPLITT Split_289_n616(net286,net169_c1,net291_c1);
SPLITT Split_297_n624(net53,net168_c1,net292_c1);
SPLITT Split_377_n704(net402,net165_c1,net293_c1);
SPLITT Split_369_n696(net382,net261_c1,net386_c1);
SPLITT Split_298_n625(net69,net175_c1,net297_c1);
SPLITT Split_378_n705(net293,net176_c1,net298_c1);
SPLITT Split_299_n626(net73,net182_c1,net303_c1);
SPLITT Split_379_n706(net165,net177_c1,net304_c1);
NOTT NOTT_140_n173(net538,net395,net136_c1);
NOTT NOTT_141_n174(net866,net403,net138_c1);
NOTT NOTT_142_n175(net808,net401,net140_c1);
NOTT NOTT_138_n165(net693,net325,net137_c1);
DFFT DFFT_184__FPB_n511(net944,net408,net410_c1);
DFFT DFFT_176__FPB_n503(net802,net409,net411_c1);
DFFT DFFT_192__FPB_n519(net690,net361,net444_c1);
DFFT DFFT_248__FPB_n575(net992,net125,net486_c1);
DFFT DFFT_168__FPB_n495(net726,net271,net489_c1);
DFFT DFFT_193__FPB_n520(net694,net444,net413_c1);
DFFT DFFT_185__FPB_n512(net752,net371,net412_c1);
DFFT DFFT_177__FPB_n504(net816,net60,net414_c1);
DFFT DFFT_249__FPB_n576(net1006,net121,net491_c1);
DFFT DFFT_169__FPB_n496(net626,net23,net493_c1);
DFFT DFFT_194__FPB_n521(net572,net223,net417_c1);
DFFT DFFT_186__FPB_n513(net758,net412,net415_c1);
DFFT DFFT_178__FPB_n505(net860,net393,net418_c1);
SPLITT Split_264_TDO(net2,net0_c1,net266_c1);
DFFT DFFT_195__FPB_n522(net912,net227,net421_c1);
DFFT DFFT_187__FPB_n514(net750,net415,net422_c1);
DFFT DFFT_179__FPB_n506(net558,net144,net423_c1);
DFFT DFFT_196__FPB_n523(net666,net146,net425_c1);
DFFT DFFT_188__FPB_n515(net560,net347,net426_c1);
DFFT DFFT_197__FPB_n524(net676,net58,net432_c1);
DFFT DFFT_189__FPB_n516(net680,net228,net430_c1);
DFFT DFFT_198__FPB_n525(net1000,net59,net436_c1);
SPLITT SplitCLK_4_251(net1001,net1006_c1,net1005_c1);
SPLITT SplitCLK_0_252(net1002,net1003_c1,net1004_c1);
SPLITT SplitCLK_0_253(net993,net1002_c1,net1001_c1);
SPLITT SplitCLK_4_254(net995,net999_c1,net1000_c1);
SPLITT SplitCLK_4_255(net996,net998_c1,net997_c1);
SPLITT SplitCLK_6_256(net994,net995_c1,net996_c1);
SPLITT SplitCLK_4_257(net977,net994_c1,net993_c1);
SPLITT SplitCLK_4_258(net987,net991_c1,net992_c1);
SPLITT SplitCLK_0_259(net988,net989_c1,net990_c1);
SPLITT SplitCLK_0_260(net979,net988_c1,net987_c1);
SPLITT SplitCLK_4_261(net981,net985_c1,net986_c1);
SPLITT SplitCLK_4_262(net982,net983_c1,net984_c1);
SPLITT SplitCLK_2_263(net980,net981_c1,net982_c1);
SPLITT SplitCLK_2_264(net978,net979_c1,net980_c1);
SPLITT SplitCLK_6_265(net945,net977_c1,net978_c1);
SPLITT SplitCLK_4_266(net971,net976_c1,net975_c1);
SPLITT SplitCLK_4_267(net972,net974_c1,net973_c1);
SPLITT SplitCLK_6_268(net963,net971_c1,net972_c1);
SPLITT SplitCLK_4_269(net965,net969_c1,net970_c1);
SPLITT SplitCLK_4_270(net966,net967_c1,net968_c1);
SPLITT SplitCLK_0_271(net964,net965_c1,net966_c1);
SPLITT SplitCLK_4_272(net947,net964_c1,net963_c1);
SPLITT SplitCLK_0_273(net957,net961_c1,net962_c1);
SPLITT SplitCLK_4_274(net958,net959_c1,net960_c1);
SPLITT SplitCLK_6_275(net949,net957_c1,net958_c1);
SPLITT SplitCLK_4_276(net951,net955_c1,net956_c1);
SPLITT SplitCLK_4_277(net952,net954_c1,net953_c1);
SPLITT SplitCLK_4_278(net950,net952_c1,net951_c1);
SPLITT SplitCLK_2_279(net948,net950_c1,net949_c1);
SPLITT SplitCLK_4_280(net946,net948_c1,net947_c1);
SPLITT SplitCLK_6_281(net883,net946_c1,net945_c1);
SPLITT SplitCLK_4_282(net939,net943_c1,net944_c1);
SPLITT SplitCLK_0_283(net940,net941_c1,net942_c1);
SPLITT SplitCLK_0_284(net931,net940_c1,net939_c1);
SPLITT SplitCLK_4_285(net933,net938_c1,net937_c1);
SPLITT SplitCLK_4_286(net934,net936_c1,net935_c1);
SPLITT SplitCLK_2_287(net932,net933_c1,net934_c1);
SPLITT SplitCLK_2_288(net915,net932_c1,net931_c1);
SPLITT SplitCLK_4_289(net925,net930_c1,net929_c1);
SPLITT SplitCLK_4_290(net926,net928_c1,net927_c1);
SPLITT SplitCLK_6_291(net917,net925_c1,net926_c1);
SPLITT SplitCLK_4_292(net919,net923_c1,net924_c1);
SPLITT SplitCLK_4_293(net920,net921_c1,net922_c1);
SPLITT SplitCLK_6_294(net918,net919_c1,net920_c1);
SPLITT SplitCLK_6_295(net916,net917_c1,net918_c1);
SPLITT SplitCLK_6_296(net885,net915_c1,net916_c1);
SPLITT SplitCLK_4_297(net909,net913_c1,net914_c1);
SPLITT SplitCLK_4_298(net910,net912_c1,net911_c1);
SPLITT SplitCLK_6_299(net901,net909_c1,net910_c1);
SPLITT SplitCLK_4_300(net903,net907_c1,net908_c1);
SPLITT SplitCLK_4_301(net904,net906_c1,net905_c1);
SPLITT SplitCLK_6_302(net902,net903_c1,net904_c1);
SPLITT SplitCLK_4_303(net887,net902_c1,net901_c1);
SPLITT SplitCLK_4_304(net895,net899_c1,net900_c1);
SPLITT SplitCLK_4_305(net896,net897_c1,net898_c1);
SPLITT SplitCLK_6_306(net889,net895_c1,net896_c1);
SPLITT SplitCLK_4_307(net892,net893_c1,net894_c1);
SPLITT SplitCLK_2_308(net890,net892_c1,net891_c1);
SPLITT SplitCLK_6_309(net888,net889_c1,net890_c1);
SPLITT SplitCLK_4_310(net886,net888_c1,net887_c1);
SPLITT SplitCLK_2_311(net884,net886_c1,net885_c1);
SPLITT SplitCLK_6_312(net759,net883_c1,net884_c1);
SPLITT SplitCLK_4_313(net877,net881_c1,net882_c1);
SPLITT SplitCLK_0_314(net878,net880_c1,net879_c1);
SPLITT SplitCLK_0_315(net869,net878_c1,net877_c1);
SPLITT SplitCLK_4_316(net871,net875_c1,net876_c1);
SPLITT SplitCLK_4_317(net872,net874_c1,net873_c1);
SPLITT SplitCLK_4_318(net870,net872_c1,net871_c1);
SPLITT SplitCLK_4_319(net853,net869_c1,net870_c1);
SPLITT SplitCLK_4_320(net863,net867_c1,net868_c1);
SPLITT SplitCLK_4_321(net864,net865_c1,net866_c1);
SPLITT SplitCLK_6_322(net855,net863_c1,net864_c1);
SPLITT SplitCLK_4_323(net857,net861_c1,net862_c1);
SPLITT SplitCLK_4_324(net858,net860_c1,net859_c1);
SPLITT SplitCLK_4_325(net856,net858_c1,net857_c1);
SPLITT SplitCLK_2_326(net854,net856_c1,net855_c1);
SPLITT SplitCLK_6_327(net823,net853_c1,net854_c1);
SPLITT SplitCLK_4_328(net847,net852_c1,net851_c1);
SPLITT SplitCLK_4_329(net848,net850_c1,net849_c1);
SPLITT SplitCLK_6_330(net839,net847_c1,net848_c1);
SPLITT SplitCLK_4_331(net841,net845_c1,net846_c1);
SPLITT SplitCLK_4_332(net842,net844_c1,net843_c1);
SPLITT SplitCLK_4_333(net840,net842_c1,net841_c1);
SPLITT SplitCLK_0_334(net825,net839_c1,net840_c1);
SPLITT SplitCLK_4_335(net833,net838_c1,net837_c1);
SPLITT SplitCLK_4_336(net834,net835_c1,net836_c1);
SPLITT SplitCLK_6_337(net827,net833_c1,net834_c1);
SPLITT SplitCLK_4_338(net830,net831_c1,net832_c1);
SPLITT SplitCLK_4_339(net828,net829_c1,net830_c1);
SPLITT SplitCLK_2_340(net826,net828_c1,net827_c1);
SPLITT SplitCLK_4_341(net824,net826_c1,net825_c1);
SPLITT SplitCLK_0_342(net761,net823_c1,net824_c1);
SPLITT SplitCLK_4_343(net817,net822_c1,net821_c1);
SPLITT SplitCLK_0_344(net818,net820_c1,net819_c1);
SPLITT SplitCLK_6_345(net809,net817_c1,net818_c1);
SPLITT SplitCLK_4_346(net811,net815_c1,net816_c1);
SPLITT SplitCLK_4_347(net812,net813_c1,net814_c1);
SPLITT SplitCLK_6_348(net810,net811_c1,net812_c1);
SPLITT SplitCLK_4_349(net793,net810_c1,net809_c1);
SPLITT SplitCLK_4_350(net803,net808_c1,net807_c1);
SPLITT SplitCLK_4_351(net804,net805_c1,net806_c1);
SPLITT SplitCLK_6_352(net795,net803_c1,net804_c1);
SPLITT SplitCLK_4_353(net797,net801_c1,net802_c1);
SPLITT SplitCLK_4_354(net798,net800_c1,net799_c1);
SPLITT SplitCLK_2_355(net796,net797_c1,net798_c1);
SPLITT SplitCLK_6_356(net794,net795_c1,net796_c1);
SPLITT SplitCLK_6_357(net763,net793_c1,net794_c1);
SPLITT SplitCLK_4_358(net787,net792_c1,net791_c1);
SPLITT SplitCLK_4_359(net788,net789_c1,net790_c1);
SPLITT SplitCLK_2_360(net779,net787_c1,net788_c1);
SPLITT SplitCLK_4_361(net781,net785_c1,net786_c1);
SPLITT SplitCLK_4_362(net782,net784_c1,net783_c1);
SPLITT SplitCLK_4_363(net780,net782_c1,net781_c1);
SPLITT SplitCLK_0_364(net765,net779_c1,net780_c1);
SPLITT SplitCLK_4_365(net773,net778_c1,net777_c1);
SPLITT SplitCLK_4_366(net774,net776_c1,net775_c1);
SPLITT SplitCLK_6_367(net767,net773_c1,net774_c1);
SPLITT SplitCLK_4_368(net770,net772_c1,net771_c1);
SPLITT SplitCLK_6_369(net768,net770_c1,net769_c1);
SPLITT SplitCLK_6_370(net766,net767_c1,net768_c1);
SPLITT SplitCLK_4_371(net764,net766_c1,net765_c1);
SPLITT SplitCLK_4_372(net762,net763_c1,net764_c1);
SPLITT SplitCLK_4_373(net760,net762_c1,net761_c1);
SPLITT SplitCLK_0_374(net503,net759_c1,net760_c1);
SPLITT SplitCLK_4_375(net753,net758_c1,net757_c1);
SPLITT SplitCLK_0_376(net754,net755_c1,net756_c1);
SPLITT SplitCLK_0_377(net745,net754_c1,net753_c1);
SPLITT SplitCLK_4_378(net747,net752_c1,net751_c1);
SPLITT SplitCLK_4_379(net748,net750_c1,net749_c1);
SPLITT SplitCLK_4_380(net746,net748_c1,net747_c1);
SPLITT SplitCLK_6_381(net729,net746_c1,net745_c1);
SPLITT SplitCLK_4_382(net739,net743_c1,net744_c1);
SPLITT SplitCLK_4_383(net740,net742_c1,net741_c1);
SPLITT SplitCLK_6_384(net731,net739_c1,net740_c1);
SPLITT SplitCLK_4_385(net733,net737_c1,net738_c1);
SPLITT SplitCLK_4_386(net734,net736_c1,net735_c1);
SPLITT SplitCLK_4_387(net732,net734_c1,net733_c1);
SPLITT SplitCLK_6_388(net730,net732_c1,net731_c1);
SPLITT SplitCLK_6_389(net697,net729_c1,net730_c1);
SPLITT SplitCLK_4_390(net723,net727_c1,net728_c1);
SPLITT SplitCLK_4_391(net724,net726_c1,net725_c1);
SPLITT SplitCLK_6_392(net715,net723_c1,net724_c1);
SPLITT SplitCLK_4_393(net717,net722_c1,net721_c1);
SPLITT SplitCLK_4_394(net718,net719_c1,net720_c1);
SPLITT SplitCLK_4_395(net716,net718_c1,net717_c1);
SPLITT SplitCLK_0_396(net699,net715_c1,net716_c1);
SPLITT SplitCLK_4_397(net709,net714_c1,net713_c1);
SPLITT SplitCLK_4_398(net710,net712_c1,net711_c1);
SPLITT SplitCLK_2_399(net701,net709_c1,net710_c1);
SPLITT SplitCLK_4_400(net703,net708_c1,net707_c1);
SPLITT SplitCLK_4_401(net704,net705_c1,net706_c1);
SPLITT SplitCLK_2_402(net702,net703_c1,net704_c1);
SPLITT SplitCLK_2_403(net700,net702_c1,net701_c1);
SPLITT SplitCLK_4_404(net698,net700_c1,net699_c1);
SPLITT SplitCLK_6_405(net635,net697_c1,net698_c1);
SPLITT SplitCLK_4_406(net691,net695_c1,net696_c1);
SPLITT SplitCLK_0_407(net692,net693_c1,net694_c1);
SPLITT SplitCLK_0_408(net683,net692_c1,net691_c1);
SPLITT SplitCLK_4_409(net685,net690_c1,net689_c1);
SPLITT SplitCLK_4_410(net686,net687_c1,net688_c1);
SPLITT SplitCLK_4_411(net684,net686_c1,net685_c1);
SPLITT SplitCLK_6_412(net667,net683_c1,net684_c1);
SPLITT SplitCLK_4_413(net677,net681_c1,net682_c1);
SPLITT SplitCLK_4_414(net678,net680_c1,net679_c1);
SPLITT SplitCLK_2_415(net669,net677_c1,net678_c1);
SPLITT SplitCLK_4_416(net671,net675_c1,net676_c1);
SPLITT SplitCLK_4_417(net672,net673_c1,net674_c1);
SPLITT SplitCLK_4_418(net670,net672_c1,net671_c1);
SPLITT SplitCLK_2_419(net668,net670_c1,net669_c1);
SPLITT SplitCLK_6_420(net637,net667_c1,net668_c1);
SPLITT SplitCLK_0_421(net661,net665_c1,net666_c1);
SPLITT SplitCLK_4_422(net662,net664_c1,net663_c1);
SPLITT SplitCLK_4_423(net653,net662_c1,net661_c1);
SPLITT SplitCLK_4_424(net655,net659_c1,net660_c1);
SPLITT SplitCLK_4_425(net656,net657_c1,net658_c1);
SPLITT SplitCLK_4_426(net654,net656_c1,net655_c1);
SPLITT SplitCLK_6_427(net639,net653_c1,net654_c1);
SPLITT SplitCLK_4_428(net647,net652_c1,net651_c1);
SPLITT SplitCLK_4_429(net648,net649_c1,net650_c1);
SPLITT SplitCLK_6_430(net641,net647_c1,net648_c1);
SPLITT SplitCLK_4_431(net644,net646_c1,net645_c1);
SPLITT SplitCLK_4_432(net642,net643_c1,net644_c1);
SPLITT SplitCLK_2_433(net640,net642_c1,net641_c1);
SPLITT SplitCLK_4_434(net638,net640_c1,net639_c1);
SPLITT SplitCLK_2_435(net636,net638_c1,net637_c1);
SPLITT SplitCLK_6_436(net511,net635_c1,net636_c1);
SPLITT SplitCLK_4_437(net629,net634_c1,net633_c1);
SPLITT SplitCLK_4_438(net630,net631_c1,net632_c1);
SPLITT SplitCLK_4_439(net621,net630_c1,net629_c1);
SPLITT SplitCLK_0_440(net623,net627_c1,net628_c1);
SPLITT SplitCLK_4_441(net624,net625_c1,net626_c1);
SPLITT SplitCLK_4_442(net622,net624_c1,net623_c1);
SPLITT SplitCLK_6_443(net605,net621_c1,net622_c1);
SPLITT SplitCLK_4_444(net615,net619_c1,net620_c1);
SPLITT SplitCLK_4_445(net616,net618_c1,net617_c1);
SPLITT SplitCLK_6_446(net607,net615_c1,net616_c1);
SPLITT SplitCLK_4_447(net609,net613_c1,net614_c1);
SPLITT SplitCLK_4_448(net610,net611_c1,net612_c1);
SPLITT SplitCLK_4_449(net608,net610_c1,net609_c1);
SPLITT SplitCLK_2_450(net606,net608_c1,net607_c1);
SPLITT SplitCLK_6_451(net575,net605_c1,net606_c1);
SPLITT SplitCLK_4_452(net599,net604_c1,net603_c1);
SPLITT SplitCLK_4_453(net600,net601_c1,net602_c1);
SPLITT SplitCLK_4_454(net591,net600_c1,net599_c1);
SPLITT SplitCLK_4_455(net593,net598_c1,net597_c1);
SPLITT SplitCLK_4_456(net594,net596_c1,net595_c1);
SPLITT SplitCLK_4_457(net592,net594_c1,net593_c1);
SPLITT SplitCLK_0_458(net577,net591_c1,net592_c1);
SPLITT SplitCLK_4_459(net585,net589_c1,net590_c1);
SPLITT SplitCLK_4_460(net586,net588_c1,net587_c1);
SPLITT SplitCLK_6_461(net579,net585_c1,net586_c1);
SPLITT SplitCLK_4_462(net582,net583_c1,net584_c1);
SPLITT SplitCLK_2_463(net580,net581_c1,net582_c1);
SPLITT SplitCLK_2_464(net578,net580_c1,net579_c1);
SPLITT SplitCLK_4_465(net576,net578_c1,net577_c1);
SPLITT SplitCLK_6_466(net513,net575_c1,net576_c1);
SPLITT SplitCLK_4_467(net569,net573_c1,net574_c1);
SPLITT SplitCLK_4_468(net570,net572_c1,net571_c1);
SPLITT SplitCLK_2_469(net561,net569_c1,net570_c1);
SPLITT SplitCLK_4_470(net563,net567_c1,net568_c1);
SPLITT SplitCLK_4_471(net564,net565_c1,net566_c1);
SPLITT SplitCLK_4_472(net562,net564_c1,net563_c1);
SPLITT SplitCLK_0_473(net545,net561_c1,net562_c1);
SPLITT SplitCLK_4_474(net555,net559_c1,net560_c1);
SPLITT SplitCLK_4_475(net556,net557_c1,net558_c1);
SPLITT SplitCLK_2_476(net547,net555_c1,net556_c1);
SPLITT SplitCLK_4_477(net549,net553_c1,net554_c1);
SPLITT SplitCLK_4_478(net550,net551_c1,net552_c1);
SPLITT SplitCLK_4_479(net548,net550_c1,net549_c1);
SPLITT SplitCLK_2_480(net546,net548_c1,net547_c1);
SPLITT SplitCLK_6_481(net515,net545_c1,net546_c1);
SPLITT SplitCLK_4_482(net539,net544_c1,net543_c1);
SPLITT SplitCLK_4_483(net540,net542_c1,net541_c1);
SPLITT SplitCLK_6_484(net531,net539_c1,net540_c1);
SPLITT SplitCLK_4_485(net533,net537_c1,net538_c1);
SPLITT SplitCLK_4_486(net534,net536_c1,net535_c1);
SPLITT SplitCLK_4_487(net532,net534_c1,net533_c1);
SPLITT SplitCLK_0_488(net517,net531_c1,net532_c1);
SPLITT SplitCLK_4_489(net525,net529_c1,net530_c1);
SPLITT SplitCLK_4_490(net526,net527_c1,net528_c1);
SPLITT SplitCLK_6_491(net519,net525_c1,net526_c1);
SPLITT SplitCLK_4_492(net522,net524_c1,net523_c1);
SPLITT SplitCLK_2_493(net520,net521_c1,net522_c1);
SPLITT SplitCLK_2_494(net518,net520_c1,net519_c1);
SPLITT SplitCLK_4_495(net516,net518_c1,net517_c1);
SPLITT SplitCLK_2_496(net514,net516_c1,net515_c1);
SPLITT SplitCLK_4_497(net512,net514_c1,net513_c1);
SPLITT SplitCLK_2_498(net504,net512_c1,net511_c1);
wire dummy0;
SPLITT SplitCLK_2_499(net769,net510_c1,dummy0);
wire dummy1;
SPLITT SplitCLK_4_500(net643,net509_c1,dummy1);
wire dummy2;
SPLITT SplitCLK_2_501(net891,net508_c1,dummy2);
wire dummy3;
SPLITT SplitCLK_2_502(net581,net507_c1,dummy3);
wire dummy4;
SPLITT SplitCLK_2_503(net521,net506_c1,dummy4);
wire dummy5;
SPLITT SplitCLK_2_504(net829,net505_c1,dummy5);
SPLITT SplitCLK_0_505(net1007,net503_c1,net504_c1);
wire dummy6;
SPLITT Split_HOLD_635(net7,dummy6,net1008_c1);
INTERCONNECT Split_264_TDO_OR2T_26_n38(net0_c1,net0);
INTERCONNECT TMS_Pad_Split_254_n581(TMS_Pad,net1);
INTERCONNECT AND2T_8_n20_Split_264_TDO(net2_c1,net2);
INTERCONNECT OR2T_9_n21_Split_265_n592(net3_c1,net3);
INTERCONNECT OR2T_18_n30_OR2T_19_n31(net4_c1,net4);
INTERCONNECT OR2T_10_n22_Split_266_n593(net5_c1,net5);
INTERCONNECT OR2T_19_n31_AND2T_22_n34(net6_c1,net6);
INTERCONNECT OR2T_11_n23_Split_HOLD_635(net7_c1,net7);
INTERCONNECT AND2T_28_n40_Split_276_n603(net8_c1,net8);
INTERCONNECT OR2T_20_n32_Split_269_n596(net9_c1,net9);
INTERCONNECT NOTT_12_n24_AND2T_134_n161(net10_c1,net10);
INTERCONNECT AND2T_4_n16_Split_256_n583(net11_c1,net11);
INTERCONNECT XOR2T_29_n41_AND2T_28_n40(net12_c1,net12);
INTERCONNECT OR2T_21_n33_AND2T_22_n34(net13_c1,net13);
INTERCONNECT OR2T_13_n25_Split_268_n595(net14_c1,net14);
INTERCONNECT NOTT_5_n17_AND2T_136_n163(net15_c1,net15);
INTERCONNECT AND2T_38_n50_Split_283_n610(net16_c1,net16);
INTERCONNECT OR2T_30_n42_Split_277_n604(net17_c1,net17);
INTERCONNECT AND2T_22_n34_AND2T_23_n35(net18_c1,net18);
INTERCONNECT OR2T_14_n26_AND2T_15_n27(net19_c1,net19);
INTERCONNECT NOTT_6_n18_Split_258_n585(net20_c1,net20);
INTERCONNECT NOTT_39_n51_AND2T_40_n52(net21_c1,net21);
INTERCONNECT AND2T_31_n43_Split_278_n605(net22_c1,net22);
INTERCONNECT AND2T_23_n35_DFFT_169__FPB_n496(net23_c1,net23);
INTERCONNECT AND2T_15_n27_AND2T_23_n35(net24_c1,net24);
INTERCONNECT AND2T_7_n19_Split_261_n588(net25_c1,net25);
INTERCONNECT AND2T_48_n60_Split_291_n618(net26_c1,net26);
INTERCONNECT AND2T_40_n52_AND2T_41_n53(net27_c1,net27);
INTERCONNECT NOTT_32_n44_AND2T_31_n43(net28_c1,net28);
INTERCONNECT AND2T_24_n36_AND2T_113_n125(net29_c1,net29);
INTERCONNECT NOTT_16_n28_AND2T_134_n161(net30_c1,net30);
INTERCONNECT NOTT_49_n61_Split_292_n619(net31_c1,net31);
INTERCONNECT AND2T_41_n53_Split_284_n611(net32_c1,net32);
INTERCONNECT AND2T_33_n45_AND2T_107_n119(net33_c1,net33);
INTERCONNECT AND2T_25_n37_OR2T_26_n38(net34_c1,net34);
INTERCONNECT AND2T_17_n29_AND2T_63_n75(net35_c1,net35);
INTERCONNECT OR2T_58_n70_OR2T_59_n71(net36_c1,net36);
INTERCONNECT AND2T_50_n62_Split_294_n621(net37_c1,net37);
INTERCONNECT NOTT_42_n54_Split_287_n614(net38_c1,net38);
INTERCONNECT AND2T_34_n46_Split_281_n608(net39_c1,net39);
INTERCONNECT OR2T_26_n38_Split_271_n598(net40_c1,net40);
INTERCONNECT OR2T_59_n71_AND2T_60_n72(net41_c1,net41);
INTERCONNECT AND2T_51_n63_OR2T_52_n64(net42_c1,net42);
INTERCONNECT OR2T_43_n55_AND2T_45_n57(net43_c1,net43);
INTERCONNECT NOTT_35_n47_AND2T_41_n53(net44_c1,net44);
INTERCONNECT AND2T_27_n39_Split_273_n600(net45_c1,net45);
INTERCONNECT OR2T_68_n80_OR2T_69_n81(net46_c1,net46);
INTERCONNECT AND2T_60_n72_OR2T_69_n81(net47_c1,net47);
INTERCONNECT OR2T_52_n64_OR2T_53_n65(net48_c1,net48);
INTERCONNECT OR2T_44_n56_AND2T_45_n57(net49_c1,net49);
INTERCONNECT OR2T_36_n48_AND2T_40_n52(net50_c1,net50);
INTERCONNECT OR2T_69_n81_OR2T_70_n82(net51_c1,net51);
INTERCONNECT AND2T_61_n73_Split_300_n627(net52_c1,net52);
INTERCONNECT OR2T_53_n65_Split_297_n624(net53_c1,net53);
INTERCONNECT AND2T_45_n57_Split_288_n615(net54_c1,net54);
INTERCONNECT AND2T_37_n49_Split_282_n609(net55_c1,net55);
INTERCONNECT OR2T_78_n90_Split_306_n633(net56_c1,net56);
INTERCONNECT OR2T_70_n82_OR2T_71_n83(net57_c1,net57);
INTERCONNECT AND2T_62_n74_DFFT_197__FPB_n524(net58_c1,net58);
INTERCONNECT AND2T_54_n66_DFFT_198__FPB_n525(net59_c1,net59);
INTERCONNECT AND2T_46_n58_DFFT_177__FPB_n504(net60_c1,net60);
INTERCONNECT OR2T_79_n91_Split_307_n634(net61_c1,net61);
INTERCONNECT OR2T_71_n83_AND2T_83_n95(net62_c1,net62);
INTERCONNECT AND2T_63_n75_Split_302_n629(net63_c1,net63);
INTERCONNECT OR2T_55_n67_AND2T_60_n72(net64_c1,net64);
INTERCONNECT AND2T_47_n59_AND2T_46_n58(net65_c1,net65);
INTERCONNECT OR2T_80_n92_Split_308_n635(net66_c1,net66);
INTERCONNECT AND2T_72_n84_Split_304_n631(net67_c1,net67);
INTERCONNECT AND2T_64_n76_AND2T_65_n77(net68_c1,net68);
INTERCONNECT AND2T_56_n68_Split_298_n625(net69_c1,net69);
INTERCONNECT OR2T_81_n93_DFFT_251__FPB_n578(net70_c1,net70);
INTERCONNECT OR2T_73_n85_OR2T_77_n89(net71_c1,net71);
INTERCONNECT AND2T_65_n77_Split_303_n630(net72_c1,net72);
INTERCONNECT AND2T_57_n69_Split_299_n626(net73_c1,net73);
INTERCONNECT OR2T_82_n94_AND2T_83_n95(net74_c1,net74);
INTERCONNECT AND2T_74_n86_OR2T_76_n88(net75_c1,net75);
INTERCONNECT OR2T_66_n78_OR2T_67_n79(net76_c1,net76);
INTERCONNECT AND2T_83_n95_Split_310_n637(net77_c1,net77);
INTERCONNECT AND2T_75_n87_Split_305_n632(net78_c1,net78);
INTERCONNECT OR2T_67_n79_OR2T_68_n80(net79_c1,net79);
INTERCONNECT AND2T_84_n96_OR2T_86_n98(net80_c1,net80);
INTERCONNECT OR2T_76_n88_OR2T_77_n89(net81_c1,net81);
INTERCONNECT AND2T_85_n97_Split_312_n639(net82_c1,net82);
INTERCONNECT OR2T_77_n89_OR2T_78_n90(net83_c1,net83);
INTERCONNECT OR2T_86_n98_Split_313_n640(net84_c1,net84);
INTERCONNECT AND2T_87_n99_DFFT_211__FPB_n538(net85_c1,net85);
INTERCONNECT AND2T_88_n100_Split_314_n641(net86_c1,net86);
INTERCONNECT AND2T_89_n101_Split_315_n642(net87_c1,net87);
INTERCONNECT AND2T_98_n110_DFFT_221__FPB_n548(net88_c1,net88);
INTERCONNECT OR2T_90_n102_OR2T_91_n103(net89_c1,net89);
INTERCONNECT AND2T_99_n111_OR2T_100_n112(net90_c1,net90);
INTERCONNECT OR2T_91_n103_OR2T_92_n104(net91_c1,net91);
INTERCONNECT OR2T_108_n120_OR2T_109_n121(net92_c1,net92);
INTERCONNECT OR2T_100_n112_OR2T_101_n113(net93_c1,net93);
INTERCONNECT OR2T_92_n104_OR2T_93_n105(net94_c1,net94);
INTERCONNECT OR2T_109_n121_DFFT_235__FPB_n562(net95_c1,net95);
INTERCONNECT OR2T_101_n113_Split_316_n643(net96_c1,net96);
INTERCONNECT OR2T_93_n105_AND2T_94_n106(net97_c1,net97);
INTERCONNECT OR2T_118_n130_AND2T_119_n131(net98_c1,net98);
INTERCONNECT AND2T_110_n122_OR2T_111_n123(net99_c1,net99);
INTERCONNECT AND2T_102_n114_AND2T_103_n115(net100_c1,net100);
INTERCONNECT AND2T_94_n106_DFFT_222__FPB_n549(net101_c1,net101);
INTERCONNECT AND2T_119_n131_Split_321_n648(net102_c1,net102);
INTERCONNECT OR2T_111_n123_OR2T_116_n128(net103_c1,net103);
INTERCONNECT AND2T_103_n115_DFFT_227__FPB_n554(net104_c1,net104);
INTERCONNECT AND2T_95_n107_AND2T_96_n108(net105_c1,net105);
INTERCONNECT OR2T_128_n140_OR2T_129_n141(net106_c1,net106);
INTERCONNECT AND2T_120_n132_AND2T_121_n133(net107_c1,net107);
INTERCONNECT AND2T_112_n124_OR2T_115_n127(net108_c1,net108);
INTERCONNECT AND2T_104_n116_Split_319_n646(net109_c1,net109);
INTERCONNECT AND2T_96_n108_OR2T_100_n112(net110_c1,net110);
INTERCONNECT OR2T_129_n141_OR2T_130_n142(net111_c1,net111);
INTERCONNECT AND2T_121_n133_DFFT_241__FPB_n568(net112_c1,net112);
INTERCONNECT AND2T_113_n125_Split_320_n647(net113_c1,net113);
INTERCONNECT OR2T_105_n117_AND2T_119_n131(net114_c1,net114);
INTERCONNECT AND2T_97_n109_AND2T_98_n110(net115_c1,net115);
INTERCONNECT OR2T_130_n142_DFFT_250__FPB_n577(net116_c1,net116);
INTERCONNECT AND2T_122_n134_Split_324_n651(net117_c1,net117);
INTERCONNECT AND2T_114_n126_OR2T_115_n127(net118_c1,net118);
INTERCONNECT AND2T_106_n118_AND2T_107_n119(net119_c1,net119);
INTERCONNECT OR2T_131_n143_AND2T_133_n145(net120_c1,net120);
INTERCONNECT AND2T_123_n135_DFFT_249__FPB_n576(net121_c1,net121);
INTERCONNECT OR2T_115_n127_OR2T_116_n128(net122_c1,net122);
INTERCONNECT AND2T_107_n119_OR2T_108_n120(net123_c1,net123);
INTERCONNECT OR2T_132_n144_AND2T_133_n145(net124_c1,net124);
INTERCONNECT AND2T_124_n136_DFFT_248__FPB_n575(net125_c1,net125);
INTERCONNECT OR2T_116_n128_OR2T_117_n129(net126_c1,net126);
INTERCONNECT AND2T_134_n161_Split_327_n654(net127_c1,net127);
INTERCONNECT AND2T_133_n145_Split_325_n652(net128_c1,net128);
INTERCONNECT AND2T_125_n137_OR2T_127_n139(net129_c1,net129);
INTERCONNECT OR2T_117_n129_DFFT_236__FPB_n563(net130_c1,net130);
INTERCONNECT AND2T_135_n162_Split_330_n657(net131_c1,net131);
INTERCONNECT OR2T_126_n138_AND2T_125_n137(net132_c1,net132);
INTERCONNECT AND2T_136_n163_Split_333_n660(net133_c1,net133);
INTERCONNECT OR2T_127_n139_OR2T_128_n140(net134_c1,net134);
INTERCONNECT AND2T_137_n164_Split_336_n663(net135_c1,net135);
INTERCONNECT NOTT_140_n173_Split_345_n672(net136_c1,net136);
INTERCONNECT NOTT_138_n165_Split_339_n666(net137_c1,net137);
INTERCONNECT NOTT_141_n174_Split_348_n675(net138_c1,net138);
INTERCONNECT OR2T_139_n166_Split_342_n669(net139_c1,net139);
INTERCONNECT NOTT_142_n175_Split_351_n678(net140_c1,net140);
INTERCONNECT Split_273_n600_Split_275_n602(net141_c1,net141);
INTERCONNECT Split_274_n601_AND2T_61_n73(net142_c1,net142);
INTERCONNECT Split_275_n602_AND2T_89_n101(net143_c1,net143);
INTERCONNECT Split_283_n610_DFFT_179__FPB_n506(net144_c1,net144);
INTERCONNECT Split_284_n611_Split_286_n613(net145_c1,net145);
INTERCONNECT Split_276_n603_DFFT_196__FPB_n523(net146_c1,net146);
INTERCONNECT Split_293_n620_DFFT_230__FPB_n557(net147_c1,net147);
INTERCONNECT Split_285_n612_AND2T_98_n110(net148_c1,net148);
INTERCONNECT Split_277_n604_OR2T_78_n90(net149_c1,net149);
INTERCONNECT Split_373_n700_DFFT_173__FPB_n500(net150_c1,net150);
INTERCONNECT Split_374_n701_Split_376_n703(net151_c1,net151);
INTERCONNECT Split_294_n621_Split_296_n623(net152_c1,net152);
INTERCONNECT Split_278_n605_Split_280_n607(net153_c1,net153);
INTERCONNECT Split_286_n613_AND2T_121_n133(net154_c1,net154);
INTERCONNECT Split_303_n630_OR2T_90_n102(net155_c1,net155);
INTERCONNECT Split_295_n622_AND2T_57_n69(net156_c1,net156);
INTERCONNECT Split_279_n606_AND2T_99_n111(net157_c1,net157);
INTERCONNECT Split_287_n614_OR2T_44_n56(net158_c1,net158);
INTERCONNECT Split_375_n702_OR2T_10_n22(net159_c1,net159);
INTERCONNECT Split_288_n615_Split_290_n617(net160_c1,net160);
INTERCONNECT Split_280_n607_AND2T_122_n134(net161_c1,net161);
INTERCONNECT Split_296_n623_AND2T_85_n97(net162_c1,net162);
INTERCONNECT Split_304_n631_OR2T_127_n139(net163_c1,net163);
INTERCONNECT Split_376_n703_DFFT_164__FPB_n491(net164_c1,net164);
INTERCONNECT Split_377_n704_Split_379_n706(net165_c1,net165);
INTERCONNECT Split_313_n640_AND2T_123_n135(net166_c1,net166);
INTERCONNECT Split_305_n632_AND2T_88_n100(net167_c1,net167);
INTERCONNECT Split_297_n624_OR2T_80_n92(net168_c1,net168);
INTERCONNECT Split_289_n616_AND2T_97_n109(net169_c1,net169);
INTERCONNECT Split_281_n608_DFFT_180__FPB_n507(net170_c1,net170);
INTERCONNECT Split_282_n609_DFFT_247__FPB_n574(net171_c1,net171);
INTERCONNECT Split_314_n641_DFFT_210__FPB_n537(net172_c1,net172);
INTERCONNECT Split_290_n617_AND2T_120_n132(net173_c1,net173);
INTERCONNECT Split_306_n633_OR2T_139_n166(net174_c1,net174);
INTERCONNECT Split_298_n625_DFFT_191__FPB_n518(net175_c1,net175);
INTERCONNECT Split_378_n705_OR2T_9_n21(net176_c1,net176);
INTERCONNECT Split_379_n706_DFFT_165__FPB_n492(net177_c1,net177);
INTERCONNECT Split_323_n650_DFFT_158__FBL_n485(net178_c1,net178);
INTERCONNECT Split_307_n634_DFFT_202__FPB_n529(net179_c1,net179);
INTERCONNECT Split_315_n642_AND2T_112_n124(net180_c1,net180);
INTERCONNECT Split_291_n618_OR2T_82_n94(net181_c1,net181);
INTERCONNECT Split_299_n626_OR2T_79_n91(net182_c1,net182);
INTERCONNECT Split_316_n643_Split_318_n645(net183_c1,net183);
INTERCONNECT Split_292_n619_Split_293_n620(net184_c1,net184);
INTERCONNECT Split_300_n627_Split_301_n628(net185_c1,net185);
INTERCONNECT Split_308_n635_Split_309_n636(net186_c1,net186);
INTERCONNECT Split_324_n651_OR2T_132_n144(net187_c1,net187);
INTERCONNECT Split_333_n660_Split_335_n662(net188_c1,net188);
INTERCONNECT Split_325_n652_Split_326_n653(net189_c1,net189);
INTERCONNECT Split_317_n644_DFFT_150__FBL_n477(net190_c1,net190);
INTERCONNECT Split_309_n636_AND2T_95_n107(net191_c1,net191);
INTERCONNECT Split_301_n628_OR2T_108_n120(net192_c1,net192);
INTERCONNECT Split_310_n637_Split_311_n638(net193_c1,net193);
INTERCONNECT Split_318_n645_DFFT_157__FBL_n484(net194_c1,net194);
INTERCONNECT Split_326_n653_DFFT_153__FBL_n480(net195_c1,net195);
INTERCONNECT Split_254_n581_Split_255_n582(net196_c1,net196);
INTERCONNECT Split_302_n629_OR2T_79_n91(net197_c1,net197);
INTERCONNECT Split_334_n661_AND2T_65_n77(net198_c1,net198);
INTERCONNECT Split_327_n654_Split_329_n656(net199_c1,net199);
INTERCONNECT Split_311_n638_DFFT_149__FBL_n476(net200_c1,net200);
INTERCONNECT Split_255_n582_DFFT_143__FPB_n185(net201_c1,net201);
INTERCONNECT Split_319_n646_OR2T_118_n130(net202_c1,net202);
INTERCONNECT Split_343_n670_AND2T_96_n108(net203_c1,net203);
INTERCONNECT Split_335_n662_AND2T_75_n87(net204_c1,net204);
INTERCONNECT Split_263_n590_AND2T_84_n96(net205_c1,net205);
INTERCONNECT Split_336_n663_Split_338_n665(net206_c1,net206);
INTERCONNECT Split_256_n583_Split_257_n584(net207_c1,net207);
INTERCONNECT Split_344_n671_DFFT_228__FPB_n555(net208_c1,net208);
INTERCONNECT Split_320_n647_AND2T_124_n136(net209_c1,net209);
INTERCONNECT Split_312_n639_AND2T_110_n122(net210_c1,net210);
INTERCONNECT Split_328_n655_AND2T_25_n37(net211_c1,net211);
INTERCONNECT Split_345_n672_Split_347_n674(net212_c1,net212);
INTERCONNECT Split_321_n648_Split_323_n650(net213_c1,net213);
INTERCONNECT Split_257_n584_DFFT_159__FPB_n486(net214_c1,net214);
INTERCONNECT Split_337_n664_NOTT_42_n54(net215_c1,net215);
INTERCONNECT Split_329_n656_AND2T_56_n68(net216_c1,net216);
INTERCONNECT Split_353_n680_OR2T_126_n138(net217_c1,net217);
INTERCONNECT Split_265_n592_DFFT_171__FPB_n498(net218_c1,net218);
INTERCONNECT Split_354_n681_Split_356_n683(net219_c1,net219);
INTERCONNECT Split_330_n657_Split_332_n659(net220_c1,net220);
INTERCONNECT Split_258_n585_Split_260_n587(net221_c1,net221);
INTERCONNECT Split_266_n593_Split_267_n594(net222_c1,net222);
INTERCONNECT Split_338_n665_DFFT_194__FPB_n521(net223_c1,net223);
INTERCONNECT Split_322_n649_DFFT_152__FBL_n479(net224_c1,net224);
INTERCONNECT Split_346_n673_OR2T_18_n30(net225_c1,net225);
INTERCONNECT Split_339_n666_Split_341_n668(net226_c1,net226);
INTERCONNECT Split_363_n690_DFFT_195__FPB_n522(net227_c1,net227);
INTERCONNECT Split_355_n682_DFFT_189__FPB_n516(net228_c1,net228);
INTERCONNECT Split_347_n674_AND2T_33_n45(net229_c1,net229);
INTERCONNECT Split_331_n658_AND2T_61_n73(net230_c1,net230);
INTERCONNECT Split_267_n594_DFFT_172__FPB_n499(net231_c1,net231);
INTERCONNECT Split_259_n586_OR2T_13_n25(net232_c1,net232);
INTERCONNECT Split_348_n675_Split_350_n677(net233_c1,net233);
INTERCONNECT Split_364_n691_DFFT_217__FPB_n544(net234_c1,net234);
INTERCONNECT Split_356_n683_DFFT_212__FPB_n539(net235_c1,net235);
INTERCONNECT Split_332_n659_AND2T_85_n97(net236_c1,net236);
INTERCONNECT Split_340_n667_DFFT_181__FPB_n508(net237_c1,net237);
INTERCONNECT Split_260_n587_AND2T_135_n162(net238_c1,net238);
INTERCONNECT Split_268_n595_OR2T_21_n33(net239_c1,net239);
INTERCONNECT Split_365_n692_Split_367_n694(net240_c1,net240);
INTERCONNECT Split_357_n684_Split_359_n686(net241_c1,net241);
INTERCONNECT Split_261_n588_Split_263_n590(net242_c1,net242);
INTERCONNECT Split_341_n668_DFFT_204__FPB_n531(net243_c1,net243);
INTERCONNECT Split_269_n596_Split_270_n597(net244_c1,net244);
INTERCONNECT Split_349_n676_AND2T_50_n62(net245_c1,net245);
INTERCONNECT Split_342_n669_Split_344_n671(net246_c1,net246);
INTERCONNECT Split_350_n677_DFFT_161__FPB_n488(net247_c1,net247);
INTERCONNECT Split_358_n685_DFFT_231__FPB_n558(net248_c1,net248);
INTERCONNECT Split_270_n597_OR2T_36_n48(net249_c1,net249);
INTERCONNECT Split_262_n589_AND2T_51_n63(net250_c1,net250);
INTERCONNECT Split_366_n693_OR2T_9_n21(net251_c1,net251);
INTERCONNECT Split_351_n678_Split_353_n680(net252_c1,net252);
INTERCONNECT Split_359_n686_DFFT_245__FPB_n572(net253_c1,net253);
INTERCONNECT Split_367_n694_DFFT_167__FPB_n494(net254_c1,net254);
INTERCONNECT Split_271_n598_Split_272_n599(net255_c1,net255);
INTERCONNECT Split_368_n695_Split_370_n697(net256_c1,net256);
INTERCONNECT Split_360_n687_Split_361_n688(net257_c1,net257);
INTERCONNECT Split_272_n599_OR2T_55_n67(net258_c1,net258);
INTERCONNECT Split_352_n679_OR2T_20_n32(net259_c1,net259);
INTERCONNECT Split_361_n688_AND2T_137_n164(net260_c1,net260);
INTERCONNECT Split_369_n696_DFFT_170__FPB_n497(net261_c1,net261);
INTERCONNECT Split_362_n689_Split_364_n691(net262_c1,net262);
INTERCONNECT Split_370_n697_DFFT_253__FPB_n580(net263_c1,net263);
INTERCONNECT Split_371_n698_Split_373_n700(net264_c1,net264);
INTERCONNECT Split_372_n699_OR2T_10_n22(net265_c1,net265);
INTERCONNECT Split_264_TDO_TDO_Pad(net266_c1,TDO_Pad);
INTERCONNECT Split_273_n600_Split_274_n601(net267_c1,net267);
INTERCONNECT Split_274_n601_AND2T_28_n40(net268_c1,net268);
INTERCONNECT Split_275_n602_AND2T_84_n96(net269_c1,net269);
INTERCONNECT Split_283_n610_NOTT_39_n51(net270_c1,net270);
INTERCONNECT Split_276_n603_DFFT_168__FPB_n495(net271_c1,net271);
INTERCONNECT Split_284_n611_Split_285_n612(net272_c1,net272);
INTERCONNECT Split_277_n604_NOTT_32_n44(net273_c1,net273);
INTERCONNECT Split_285_n612_AND2T_46_n58(net274_c1,net274);
INTERCONNECT Split_293_n620_DFFT_207__FPB_n534(net275_c1,net275);
INTERCONNECT Split_373_n700_NOTT_16_n28(net276_c1,net276);
INTERCONNECT Split_278_n605_Split_279_n606(net277_c1,net277);
INTERCONNECT Split_286_n613_AND2T_103_n115(net278_c1,net278);
INTERCONNECT Split_294_n621_Split_295_n622(net279_c1,net279);
INTERCONNECT Split_374_n701_Split_375_n702(net280_c1,net280);
INTERCONNECT Split_279_n606_AND2T_48_n60(net281_c1,net281);
INTERCONNECT Split_287_n614_OR2T_43_n55(net282_c1,net282);
INTERCONNECT Split_295_n622_AND2T_51_n63(net283_c1,net283);
INTERCONNECT Split_375_n702_AND2T_4_n16(net284_c1,net284);
INTERCONNECT Split_303_n630_OR2T_66_n78(net285_c1,net285);
INTERCONNECT Split_288_n615_Split_289_n616(net286_c1,net286);
INTERCONNECT Split_296_n623_AND2T_75_n87(net287_c1,net287);
INTERCONNECT Split_376_n703_NOTT_12_n24(net288_c1,net288);
INTERCONNECT Split_280_n607_AND2T_104_n116(net289_c1,net289);
INTERCONNECT Split_304_n631_OR2T_73_n85(net290_c1,net290);
INTERCONNECT Split_289_n616_AND2T_47_n59(net291_c1,net291);
INTERCONNECT Split_297_n624_AND2T_54_n66(net292_c1,net292);
INTERCONNECT Split_377_n704_Split_378_n705(net293_c1,net293);
INTERCONNECT Split_281_n608_NOTT_35_n47(net294_c1,net294);
INTERCONNECT Split_305_n632_OR2T_76_n88(net295_c1,net295);
INTERCONNECT Split_313_n640_AND2T_87_n99(net296_c1,net296);
INTERCONNECT Split_298_n625_OR2T_73_n85(net297_c1,net297);
INTERCONNECT Split_378_n705_NOTT_5_n17(net298_c1,net298);
INTERCONNECT Split_282_n609_DFFT_208__FPB_n535(net299_c1,net299);
INTERCONNECT Split_290_n617_AND2T_102_n114(net300_c1,net300);
INTERCONNECT Split_306_n633_OR2T_81_n93(net301_c1,net301);
INTERCONNECT Split_314_n641_OR2T_128_n140(net302_c1,net302);
INTERCONNECT Split_299_n626_OR2T_58_n70(net303_c1,net303);
INTERCONNECT Split_379_n706_DFFT_160__FPB_n487(net304_c1,net304);
INTERCONNECT Split_291_n618_OR2T_71_n83(net305_c1,net305);
INTERCONNECT Split_307_n634_OR2T_111_n123(net306_c1,net306);
INTERCONNECT Split_315_n642_OR2T_90_n102(net307_c1,net307);
INTERCONNECT Split_323_n650_DFFT_154__FBL_n481(net308_c1,net308);
INTERCONNECT Split_292_n619_DFFT_234__FPB_n561(net309_c1,net309);
INTERCONNECT Split_308_n635_OR2T_139_n166(net310_c1,net310);
INTERCONNECT Split_316_n643_Split_317_n644(net311_c1,net311);
INTERCONNECT Split_324_n651_OR2T_131_n143(net312_c1,net312);
INTERCONNECT Split_300_n627_DFFT_209__FPB_n536(net313_c1,net313);
INTERCONNECT Split_309_n636_OR2T_81_n93(net314_c1,net314);
INTERCONNECT Split_317_n644_DFFT_146__FBL_n473(net315_c1,net315);
INTERCONNECT Split_325_n652_DFFT_155__FBL_n482(net316_c1,net316);
INTERCONNECT Split_333_n660_Split_334_n661(net317_c1,net317);
INTERCONNECT Split_301_n628_AND2T_62_n74(net318_c1,net318);
INTERCONNECT Split_254_n581_DFFT_144__FPB_n186(net319_c1,net319);
INTERCONNECT Split_318_n645_DFFT_151__FBL_n478(net320_c1,net320);
INTERCONNECT Split_326_n653_DFFT_148__FBL_n475(net321_c1,net321);
INTERCONNECT Split_334_n661_AND2T_34_n46(net322_c1,net322);
INTERCONNECT Split_302_n629_OR2T_66_n78(net323_c1,net323);
INTERCONNECT Split_310_n637_DFFT_156__FBL_n483(net324_c1,net324);
INTERCONNECT Split_255_n582_NOTT_138_n165(net325_c1,net325);
INTERCONNECT Split_263_n590_AND2T_56_n68(net326_c1,net326);
INTERCONNECT Split_319_n646_OR2T_105_n117(net327_c1,net327);
INTERCONNECT Split_327_n654_Split_328_n655(net328_c1,net328);
INTERCONNECT Split_335_n662_AND2T_72_n84(net329_c1,net329);
INTERCONNECT Split_343_n670_AND2T_94_n106(net330_c1,net330);
INTERCONNECT Split_311_n638_DFFT_145__FBL_n472(net331_c1,net331);
INTERCONNECT Split_256_n583_DFFT_233__FPB_n560(net332_c1,net332);
INTERCONNECT Split_328_n655_OR2T_19_n31(net333_c1,net333);
INTERCONNECT Split_336_n663_Split_337_n664(net334_c1,net334);
INTERCONNECT Split_344_n671_DFFT_203__FPB_n530(net335_c1,net335);
INTERCONNECT Split_312_n639_OR2T_86_n98(net336_c1,net336);
INTERCONNECT Split_320_n647_AND2T_114_n126(net337_c1,net337);
INTERCONNECT Split_257_n584_AND2T_38_n50(net338_c1,net338);
INTERCONNECT Split_265_n592_OR2T_11_n23(net339_c1,net339);
INTERCONNECT Split_329_n656_AND2T_34_n46(net340_c1,net340);
INTERCONNECT Split_337_n664_AND2T_38_n50(net341_c1,net341);
INTERCONNECT Split_345_n672_Split_346_n673(net342_c1,net342);
INTERCONNECT Split_353_n680_AND2T_27_n39(net343_c1,net343);
INTERCONNECT Split_321_n648_Split_322_n649(net344_c1,net344);
INTERCONNECT Split_258_n585_Split_259_n586(net345_c1,net345);
INTERCONNECT Split_266_n593_DFFT_201__FPB_n528(net346_c1,net346);
INTERCONNECT Split_338_n665_DFFT_188__FPB_n515(net347_c1,net347);
INTERCONNECT Split_346_n673_AND2T_7_n19(net348_c1,net348);
INTERCONNECT Split_354_n681_Split_355_n682(net349_c1,net349);
INTERCONNECT Split_322_n649_DFFT_147__FBL_n474(net350_c1,net350);
INTERCONNECT Split_330_n657_Split_331_n658(net351_c1,net351);
INTERCONNECT Split_259_n586_AND2T_7_n19(net352_c1,net352);
INTERCONNECT Split_267_n594_OR2T_11_n23(net353_c1,net353);
INTERCONNECT Split_339_n666_Split_340_n667(net354_c1,net354);
INTERCONNECT Split_347_n674_XOR2T_29_n41(net355_c1,net355);
INTERCONNECT Split_355_n682_NOTT_49_n61(net356_c1,net356);
INTERCONNECT Split_363_n690_DFFT_166__FPB_n493(net357_c1,net357);
INTERCONNECT Split_331_n658_AND2T_25_n37(net358_c1,net358);
INTERCONNECT Split_268_n595_OR2T_14_n26(net359_c1,net359);
INTERCONNECT Split_348_n675_Split_349_n676(net360_c1,net360);
INTERCONNECT Split_356_n683_DFFT_192__FPB_n519(net361_c1,net361);
INTERCONNECT Split_364_n691_DFFT_199__FPB_n526(net362_c1,net362);
INTERCONNECT Split_260_n587_AND2T_24_n36(net363_c1,net363);
INTERCONNECT Split_332_n659_AND2T_74_n86(net364_c1,net364);
INTERCONNECT Split_340_n667_AND2T_64_n76(net365_c1,net365);
INTERCONNECT Split_269_n596_OR2T_43_n55(net366_c1,net366);
INTERCONNECT Split_349_n676_AND2T_17_n29(net367_c1,net367);
INTERCONNECT Split_357_n684_Split_358_n685(net368_c1,net368);
INTERCONNECT Split_365_n692_Split_366_n693(net369_c1,net369);
INTERCONNECT Split_261_n588_Split_262_n589(net370_c1,net370);
INTERCONNECT Split_341_n668_DFFT_185__FPB_n512(net371_c1,net371);
INTERCONNECT Split_358_n685_AND2T_106_n118(net372_c1,net372);
INTERCONNECT Split_366_n693_NOTT_6_n18(net373_c1,net373);
INTERCONNECT Split_262_n589_AND2T_8_n20(net374_c1,net374);
INTERCONNECT Split_270_n597_OR2T_21_n33(net375_c1,net375);
INTERCONNECT Split_342_n669_Split_343_n670(net376_c1,net376);
INTERCONNECT Split_350_n677_OR2T_126_n138(net377_c1,net377);
INTERCONNECT Split_359_n686_DFFT_242__FPB_n569(net378_c1,net378);
INTERCONNECT Split_367_n694_DFFT_163__FPB_n490(net379_c1,net379);
INTERCONNECT Split_271_n598_OR2T_109_n121(net380_c1,net380);
INTERCONNECT Split_351_n678_Split_352_n679(net381_c1,net381);
INTERCONNECT Split_368_n695_Split_369_n696(net382_c1,net382);
INTERCONNECT Split_272_n599_OR2T_30_n42(net383_c1,net383);
INTERCONNECT Split_352_n679_AND2T_17_n29(net384_c1,net384);
INTERCONNECT Split_360_n687_DFFT_223__FPB_n550(net385_c1,net385);
INTERCONNECT Split_369_n696_AND2T_37_n49(net386_c1,net386);
INTERCONNECT Split_361_n688_AND2T_37_n49(net387_c1,net387);
INTERCONNECT Split_362_n689_Split_363_n690(net388_c1,net388);
INTERCONNECT Split_370_n697_DFFT_237__FPB_n564(net389_c1,net389);
INTERCONNECT Split_371_n698_Split_372_n699(net390_c1,net390);
INTERCONNECT Split_372_n699_AND2T_4_n16(net391_c1,net391);
INTERCONNECT DFFT_153__FBL_n480_Split_365_n692(net392_c1,net392);
INTERCONNECT DFFT_145__FBL_n472_DFFT_178__FPB_n505(net393_c1,net393);
INTERCONNECT DFFT_146__FBL_n473_DFFT_229__FPB_n556(net394_c1,net394);
INTERCONNECT DFFT_154__FBL_n481_NOTT_140_n173(net395_c1,net395);
INTERCONNECT DFFT_155__FBL_n482_Split_368_n695(net396_c1,net396);
INTERCONNECT DFFT_147__FBL_n474_Split_360_n687(net397_c1,net397);
INTERCONNECT DFFT_156__FBL_n483_Split_371_n698(net398_c1,net398);
INTERCONNECT DFFT_148__FBL_n475_AND2T_137_n164(net399_c1,net399);
INTERCONNECT DFFT_157__FBL_n484_Split_374_n701(net400_c1,net400);
INTERCONNECT DFFT_149__FBL_n476_NOTT_142_n175(net401_c1,net401);
INTERCONNECT DFFT_158__FBL_n485_Split_377_n704(net402_c1,net402);
INTERCONNECT DFFT_150__FBL_n477_NOTT_141_n174(net403_c1,net403);
INTERCONNECT DFFT_151__FBL_n478_Split_362_n689(net404_c1,net404);
INTERCONNECT DFFT_152__FBL_n479_DFFT_252__FPB_n579(net405_c1,net405);
INTERCONNECT DFFT_173__FPB_n500_DFFT_174__FPB_n501(net406_c1,net406);
INTERCONNECT DFFT_174__FPB_n501_DFFT_175__FPB_n502(net407_c1,net407);
INTERCONNECT DFFT_183__FPB_n510_DFFT_184__FPB_n511(net408_c1,net408);
INTERCONNECT DFFT_175__FPB_n502_DFFT_176__FPB_n503(net409_c1,net409);
INTERCONNECT DFFT_184__FPB_n511_AND2T_54_n66(net410_c1,net410);
INTERCONNECT DFFT_176__FPB_n503_AND2T_47_n59(net411_c1,net411);
INTERCONNECT DFFT_185__FPB_n512_DFFT_186__FPB_n513(net412_c1,net412);
INTERCONNECT DFFT_193__FPB_n520_AND2T_62_n74(net413_c1,net413);
INTERCONNECT DFFT_177__FPB_n504_AND2T_48_n60(net414_c1,net414);
INTERCONNECT DFFT_186__FPB_n513_DFFT_187__FPB_n514(net415_c1,net415);
INTERCONNECT DFFT_143__FPB_n185_Split_354_n681(net416_c1,net416);
INTERCONNECT DFFT_194__FPB_n521_AND2T_63_n75(net417_c1,net417);
INTERCONNECT DFFT_178__FPB_n505_AND2T_50_n62(net418_c1,net418);
INTERCONNECT DFFT_144__FPB_n186_Split_357_n684(net419_c1,net419);
INTERCONNECT DFFT_203__FPB_n530_OR2T_82_n94(net420_c1,net420);
INTERCONNECT DFFT_195__FPB_n522_AND2T_64_n76(net421_c1,net421);
INTERCONNECT DFFT_187__FPB_n514_OR2T_55_n67(net422_c1,net422);
INTERCONNECT DFFT_179__FPB_n506_OR2T_52_n64(net423_c1,net423);
INTERCONNECT DFFT_204__FPB_n531_DFFT_205__FPB_n532(net424_c1,net424);
INTERCONNECT DFFT_196__FPB_n523_OR2T_67_n79(net425_c1,net425);
INTERCONNECT DFFT_188__FPB_n515_AND2T_57_n69(net426_c1,net426);
INTERCONNECT DFFT_180__FPB_n507_OR2T_53_n65(net427_c1,net427);
INTERCONNECT DFFT_213__FPB_n540_DFFT_214__FPB_n541(net428_c1,net428);
INTERCONNECT DFFT_205__FPB_n532_DFFT_206__FPB_n533(net429_c1,net429);
INTERCONNECT DFFT_189__FPB_n516_DFFT_190__FPB_n517(net430_c1,net430);
INTERCONNECT DFFT_181__FPB_n508_DFFT_182__FPB_n509(net431_c1,net431);
INTERCONNECT DFFT_197__FPB_n524_OR2T_68_n80(net432_c1,net432);
INTERCONNECT DFFT_214__FPB_n541_DFFT_215__FPB_n542(net433_c1,net433);
INTERCONNECT DFFT_182__FPB_n509_DFFT_183__FPB_n510(net434_c1,net434);
INTERCONNECT DFFT_206__FPB_n533_AND2T_87_n99(net435_c1,net435);
INTERCONNECT DFFT_198__FPB_n525_OR2T_70_n82(net436_c1,net436);
INTERCONNECT DFFT_190__FPB_n517_OR2T_58_n70(net437_c1,net437);
INTERCONNECT DFFT_223__FPB_n550_DFFT_224__FPB_n551(net438_c1,net438);
INTERCONNECT DFFT_215__FPB_n542_DFFT_216__FPB_n543(net439_c1,net439);
INTERCONNECT DFFT_199__FPB_n526_DFFT_200__FPB_n527(net440_c1,net440);
INTERCONNECT DFFT_207__FPB_n534_AND2T_88_n100(net441_c1,net441);
INTERCONNECT DFFT_191__FPB_n518_OR2T_59_n71(net442_c1,net442);
INTERCONNECT DFFT_224__FPB_n551_DFFT_225__FPB_n552(net443_c1,net443);
INTERCONNECT DFFT_192__FPB_n519_DFFT_193__FPB_n520(net444_c1,net444);
INTERCONNECT DFFT_216__FPB_n543_AND2T_95_n107(net445_c1,net445);
INTERCONNECT DFFT_208__FPB_n535_AND2T_89_n101(net446_c1,net446);
INTERCONNECT DFFT_200__FPB_n527_AND2T_72_n84(net447_c1,net447);
INTERCONNECT DFFT_225__FPB_n552_DFFT_226__FPB_n553(net448_c1,net448);
INTERCONNECT DFFT_217__FPB_n544_DFFT_218__FPB_n545(net449_c1,net449);
INTERCONNECT DFFT_233__FPB_n560_AND2T_113_n125(net450_c1,net450);
INTERCONNECT DFFT_209__FPB_n536_OR2T_91_n103(net451_c1,net451);
INTERCONNECT DFFT_201__FPB_n528_AND2T_74_n86(net452_c1,net452);
INTERCONNECT DFFT_218__FPB_n545_DFFT_219__FPB_n546(net453_c1,net453);
INTERCONNECT DFFT_234__FPB_n561_AND2T_114_n126(net454_c1,net454);
INTERCONNECT DFFT_226__FPB_n553_AND2T_102_n114(net455_c1,net455);
INTERCONNECT DFFT_210__FPB_n537_OR2T_92_n104(net456_c1,net456);
INTERCONNECT DFFT_202__FPB_n529_OR2T_80_n92(net457_c1,net457);
INTERCONNECT DFFT_243__FPB_n570_DFFT_244__FPB_n571(net458_c1,net458);
INTERCONNECT DFFT_219__FPB_n546_DFFT_220__FPB_n547(net459_c1,net459);
INTERCONNECT DFFT_235__FPB_n562_OR2T_117_n129(net460_c1,net460);
INTERCONNECT DFFT_227__FPB_n554_AND2T_104_n116(net461_c1,net461);
INTERCONNECT DFFT_211__FPB_n538_OR2T_93_n105(net462_c1,net462);
INTERCONNECT DFFT_163__FPB_n490_OR2T_18_n30(net463_c1,net463);
INTERCONNECT DFFT_212__FPB_n539_DFFT_213__FPB_n540(net464_c1,net464);
INTERCONNECT DFFT_244__FPB_n571_AND2T_123_n135(net465_c1,net465);
INTERCONNECT DFFT_236__FPB_n563_OR2T_118_n130(net466_c1,net466);
INTERCONNECT DFFT_228__FPB_n555_OR2T_105_n117(net467_c1,net467);
INTERCONNECT DFFT_220__FPB_n547_AND2T_97_n109(net468_c1,net468);
INTERCONNECT DFFT_164__FPB_n491_OR2T_20_n32(net469_c1,net469);
INTERCONNECT DFFT_245__FPB_n572_DFFT_246__FPB_n573(net470_c1,net470);
INTERCONNECT DFFT_237__FPB_n564_DFFT_238__FPB_n565(net471_c1,net471);
INTERCONNECT DFFT_253__FPB_n580_AND2T_136_n163(net472_c1,net472);
INTERCONNECT DFFT_229__FPB_n556_AND2T_106_n118(net473_c1,net473);
INTERCONNECT DFFT_221__FPB_n548_AND2T_99_n111(net474_c1,net474);
INTERCONNECT DFFT_165__FPB_n492_AND2T_24_n36(net475_c1,net475);
INTERCONNECT DFFT_238__FPB_n565_DFFT_239__FPB_n566(net476_c1,net476);
INTERCONNECT DFFT_246__FPB_n573_AND2T_124_n136(net477_c1,net477);
INTERCONNECT DFFT_230__FPB_n557_AND2T_110_n122(net478_c1,net478);
INTERCONNECT DFFT_222__FPB_n549_OR2T_101_n113(net479_c1,net479);
INTERCONNECT DFFT_166__FPB_n493_AND2T_27_n39(net480_c1,net480);
INTERCONNECT DFFT_239__FPB_n566_DFFT_240__FPB_n567(net481_c1,net481);
INTERCONNECT DFFT_231__FPB_n558_DFFT_232__FPB_n559(net482_c1,net482);
INTERCONNECT DFFT_247__FPB_n574_AND2T_125_n137(net483_c1,net483);
INTERCONNECT DFFT_167__FPB_n494_XOR2T_29_n41(net484_c1,net484);
INTERCONNECT DFFT_159__FPB_n486_AND2T_8_n20(net485_c1,net485);
INTERCONNECT DFFT_248__FPB_n575_OR2T_129_n141(net486_c1,net486);
INTERCONNECT DFFT_240__FPB_n567_AND2T_120_n132(net487_c1,net487);
INTERCONNECT DFFT_232__FPB_n559_AND2T_112_n124(net488_c1,net488);
INTERCONNECT DFFT_168__FPB_n495_OR2T_30_n42(net489_c1,net489);
INTERCONNECT DFFT_160__FPB_n487_OR2T_13_n25(net490_c1,net490);
INTERCONNECT DFFT_249__FPB_n576_OR2T_130_n142(net491_c1,net491);
INTERCONNECT DFFT_241__FPB_n568_AND2T_122_n134(net492_c1,net492);
INTERCONNECT DFFT_169__FPB_n496_AND2T_31_n43(net493_c1,net493);
INTERCONNECT DFFT_161__FPB_n488_OR2T_14_n26(net494_c1,net494);
INTERCONNECT DFFT_242__FPB_n569_DFFT_243__FPB_n570(net495_c1,net495);
INTERCONNECT DFFT_250__FPB_n577_OR2T_131_n143(net496_c1,net496);
INTERCONNECT DFFT_170__FPB_n497_AND2T_33_n45(net497_c1,net497);
INTERCONNECT DFFT_162__FPB_n489_AND2T_15_n27(net498_c1,net498);
INTERCONNECT DFFT_251__FPB_n578_OR2T_132_n144(net499_c1,net499);
INTERCONNECT DFFT_171__FPB_n498_OR2T_36_n48(net500_c1,net500);
INTERCONNECT DFFT_252__FPB_n579_AND2T_135_n162(net501_c1,net501);
INTERCONNECT DFFT_172__FPB_n499_OR2T_44_n56(net502_c1,net502);
INTERCONNECT SplitCLK_0_505_SplitCLK_0_374(net503_c1,net503);
INTERCONNECT SplitCLK_0_505_SplitCLK_2_498(net504_c1,net504);
INTERCONNECT SplitCLK_2_504_DFFT_167__FPB_n494(net505_c1,net505);
INTERCONNECT SplitCLK_2_503_DFFT_158__FBL_n485(net506_c1,net506);
INTERCONNECT SplitCLK_2_502_DFFT_152__FBL_n479(net507_c1,net507);
INTERCONNECT SplitCLK_2_501_AND2T_72_n84(net508_c1,net508);
INTERCONNECT SplitCLK_4_500_AND2T_8_n20(net509_c1,net509);
INTERCONNECT SplitCLK_2_499_AND2T_136_n163(net510_c1,net510);
INTERCONNECT SplitCLK_2_498_SplitCLK_6_436(net511_c1,net511);
INTERCONNECT SplitCLK_2_498_SplitCLK_4_497(net512_c1,net512);
INTERCONNECT SplitCLK_4_497_SplitCLK_6_466(net513_c1,net513);
INTERCONNECT SplitCLK_4_497_SplitCLK_2_496(net514_c1,net514);
INTERCONNECT SplitCLK_2_496_SplitCLK_6_481(net515_c1,net515);
INTERCONNECT SplitCLK_2_496_SplitCLK_4_495(net516_c1,net516);
INTERCONNECT SplitCLK_4_495_SplitCLK_0_488(net517_c1,net517);
INTERCONNECT SplitCLK_4_495_SplitCLK_2_494(net518_c1,net518);
INTERCONNECT SplitCLK_2_494_SplitCLK_6_491(net519_c1,net519);
INTERCONNECT SplitCLK_2_494_SplitCLK_2_493(net520_c1,net520);
INTERCONNECT SplitCLK_2_493_SplitCLK_2_503(net521_c1,net521);
INTERCONNECT SplitCLK_2_493_SplitCLK_4_492(net522_c1,net522);
INTERCONNECT SplitCLK_4_492_NOTT_5_n17(net523_c1,net523);
INTERCONNECT SplitCLK_4_492_DFFT_165__FPB_n492(net524_c1,net524);
INTERCONNECT SplitCLK_6_491_SplitCLK_4_489(net525_c1,net525);
INTERCONNECT SplitCLK_6_491_SplitCLK_4_490(net526_c1,net526);
INTERCONNECT SplitCLK_4_490_NOTT_42_n54(net527_c1,net527);
INTERCONNECT SplitCLK_4_490_DFFT_171__FPB_n498(net528_c1,net528);
INTERCONNECT SplitCLK_4_489_AND2T_24_n36(net529_c1,net529);
INTERCONNECT SplitCLK_4_489_OR2T_11_n23(net530_c1,net530);
INTERCONNECT SplitCLK_0_488_SplitCLK_6_484(net531_c1,net531);
INTERCONNECT SplitCLK_0_488_SplitCLK_4_487(net532_c1,net532);
INTERCONNECT SplitCLK_4_487_SplitCLK_4_485(net533_c1,net533);
INTERCONNECT SplitCLK_4_487_SplitCLK_4_486(net534_c1,net534);
INTERCONNECT SplitCLK_4_486_OR2T_9_n21(net535_c1,net535);
INTERCONNECT SplitCLK_4_486_DFFT_160__FPB_n487(net536_c1,net536);
INTERCONNECT SplitCLK_4_485_DFFT_154__FBL_n481(net537_c1,net537);
INTERCONNECT SplitCLK_4_485_NOTT_140_n173(net538_c1,net538);
INTERCONNECT SplitCLK_6_484_SplitCLK_4_482(net539_c1,net539);
INTERCONNECT SplitCLK_6_484_SplitCLK_4_483(net540_c1,net540);
INTERCONNECT SplitCLK_4_483_OR2T_13_n25(net541_c1,net541);
INTERCONNECT SplitCLK_4_483_DFFT_162__FPB_n489(net542_c1,net542);
INTERCONNECT SplitCLK_4_482_AND2T_7_n19(net543_c1,net543);
INTERCONNECT SplitCLK_4_482_OR2T_43_n55(net544_c1,net544);
INTERCONNECT SplitCLK_6_481_SplitCLK_0_473(net545_c1,net545);
INTERCONNECT SplitCLK_6_481_SplitCLK_2_480(net546_c1,net546);
INTERCONNECT SplitCLK_2_480_SplitCLK_2_476(net547_c1,net547);
INTERCONNECT SplitCLK_2_480_SplitCLK_4_479(net548_c1,net548);
INTERCONNECT SplitCLK_4_479_SplitCLK_4_477(net549_c1,net549);
INTERCONNECT SplitCLK_4_479_SplitCLK_4_478(net550_c1,net550);
INTERCONNECT SplitCLK_4_478_AND2T_38_n50(net551_c1,net551);
INTERCONNECT SplitCLK_4_478_DFFT_233__FPB_n560(net552_c1,net552);
INTERCONNECT SplitCLK_4_477_OR2T_44_n56(net553_c1,net553);
INTERCONNECT SplitCLK_4_477_NOTT_39_n51(net554_c1,net554);
INTERCONNECT SplitCLK_2_476_SplitCLK_4_474(net555_c1,net555);
INTERCONNECT SplitCLK_2_476_SplitCLK_4_475(net556_c1,net556);
INTERCONNECT SplitCLK_4_475_DFFT_159__FPB_n486(net557_c1,net557);
INTERCONNECT SplitCLK_4_475_DFFT_179__FPB_n506(net558_c1,net558);
INTERCONNECT SplitCLK_4_474_OR2T_52_n64(net559_c1,net559);
INTERCONNECT SplitCLK_4_474_DFFT_188__FPB_n515(net560_c1,net560);
INTERCONNECT SplitCLK_0_473_SplitCLK_2_469(net561_c1,net561);
INTERCONNECT SplitCLK_0_473_SplitCLK_4_472(net562_c1,net562);
INTERCONNECT SplitCLK_4_472_SplitCLK_4_470(net563_c1,net563);
INTERCONNECT SplitCLK_4_472_SplitCLK_4_471(net564_c1,net564);
INTERCONNECT SplitCLK_4_471_AND2T_113_n125(net565_c1,net565);
INTERCONNECT SplitCLK_4_471_DFFT_172__FPB_n499(net566_c1,net566);
INTERCONNECT SplitCLK_4_470_AND2T_4_n16(net567_c1,net567);
INTERCONNECT SplitCLK_4_470_AND2T_40_n52(net568_c1,net568);
INTERCONNECT SplitCLK_2_469_SplitCLK_4_467(net569_c1,net569);
INTERCONNECT SplitCLK_2_469_SplitCLK_4_468(net570_c1,net570);
INTERCONNECT SplitCLK_4_468_AND2T_57_n69(net571_c1,net571);
INTERCONNECT SplitCLK_4_468_DFFT_194__FPB_n521(net572_c1,net572);
INTERCONNECT SplitCLK_4_467_AND2T_63_n75(net573_c1,net573);
INTERCONNECT SplitCLK_4_467_OR2T_10_n22(net574_c1,net574);
INTERCONNECT SplitCLK_6_466_SplitCLK_6_451(net575_c1,net575);
INTERCONNECT SplitCLK_6_466_SplitCLK_4_465(net576_c1,net576);
INTERCONNECT SplitCLK_4_465_SplitCLK_0_458(net577_c1,net577);
INTERCONNECT SplitCLK_4_465_SplitCLK_2_464(net578_c1,net578);
INTERCONNECT SplitCLK_2_464_SplitCLK_6_461(net579_c1,net579);
INTERCONNECT SplitCLK_2_464_SplitCLK_2_463(net580_c1,net580);
INTERCONNECT SplitCLK_2_463_SplitCLK_2_502(net581_c1,net581);
INTERCONNECT SplitCLK_2_463_SplitCLK_4_462(net582_c1,net582);
INTERCONNECT SplitCLK_4_462_NOTT_6_n18(net583_c1,net583);
INTERCONNECT SplitCLK_4_462_DFFT_147__FBL_n474(net584_c1,net584);
INTERCONNECT SplitCLK_6_461_SplitCLK_4_459(net585_c1,net585);
INTERCONNECT SplitCLK_6_461_SplitCLK_4_460(net586_c1,net586);
INTERCONNECT SplitCLK_4_460_AND2T_135_n162(net587_c1,net587);
INTERCONNECT SplitCLK_4_460_AND2T_45_n57(net588_c1,net588);
INTERCONNECT SplitCLK_4_459_OR2T_21_n33(net589_c1,net589);
INTERCONNECT SplitCLK_4_459_OR2T_14_n26(net590_c1,net590);
INTERCONNECT SplitCLK_0_458_SplitCLK_4_454(net591_c1,net591);
INTERCONNECT SplitCLK_0_458_SplitCLK_4_457(net592_c1,net592);
INTERCONNECT SplitCLK_4_457_SplitCLK_4_455(net593_c1,net593);
INTERCONNECT SplitCLK_4_457_SplitCLK_4_456(net594_c1,net594);
INTERCONNECT SplitCLK_4_456_DFFT_153__FBL_n480(net595_c1,net595);
INTERCONNECT SplitCLK_4_456_DFFT_252__FPB_n579(net596_c1,net596);
INTERCONNECT SplitCLK_4_455_AND2T_15_n27(net597_c1,net597);
INTERCONNECT SplitCLK_4_455_DFFT_148__FBL_n475(net598_c1,net598);
INTERCONNECT SplitCLK_4_454_SplitCLK_4_452(net599_c1,net599);
INTERCONNECT SplitCLK_4_454_SplitCLK_4_453(net600_c1,net600);
INTERCONNECT SplitCLK_4_453_AND2T_119_n131(net601_c1,net601);
INTERCONNECT SplitCLK_4_453_AND2T_23_n35(net602_c1,net602);
INTERCONNECT SplitCLK_4_452_AND2T_22_n34(net603_c1,net603);
INTERCONNECT SplitCLK_4_452_OR2T_118_n130(net604_c1,net604);
INTERCONNECT SplitCLK_6_451_SplitCLK_6_443(net605_c1,net605);
INTERCONNECT SplitCLK_6_451_SplitCLK_2_450(net606_c1,net606);
INTERCONNECT SplitCLK_2_450_SplitCLK_6_446(net607_c1,net607);
INTERCONNECT SplitCLK_2_450_SplitCLK_4_449(net608_c1,net608);
INTERCONNECT SplitCLK_4_449_SplitCLK_4_447(net609_c1,net609);
INTERCONNECT SplitCLK_4_449_SplitCLK_4_448(net610_c1,net610);
INTERCONNECT SplitCLK_4_448_AND2T_41_n53(net611_c1,net611);
INTERCONNECT SplitCLK_4_448_OR2T_36_n48(net612_c1,net612);
INTERCONNECT SplitCLK_4_447_NOTT_35_n47(net613_c1,net613);
INTERCONNECT SplitCLK_4_447_DFFT_161__FPB_n488(net614_c1,net614);
INTERCONNECT SplitCLK_6_446_SplitCLK_4_444(net615_c1,net615);
INTERCONNECT SplitCLK_6_446_SplitCLK_4_445(net616_c1,net616);
INTERCONNECT SplitCLK_4_445_OR2T_20_n32(net617_c1,net617);
INTERCONNECT SplitCLK_4_445_DFFT_201__FPB_n528(net618_c1,net618);
INTERCONNECT SplitCLK_4_444_DFFT_180__FPB_n507(net619_c1,net619);
INTERCONNECT SplitCLK_4_444_DFFT_164__FPB_n491(net620_c1,net620);
INTERCONNECT SplitCLK_6_443_SplitCLK_4_439(net621_c1,net621);
INTERCONNECT SplitCLK_6_443_SplitCLK_4_442(net622_c1,net622);
INTERCONNECT SplitCLK_4_442_SplitCLK_0_440(net623_c1,net623);
INTERCONNECT SplitCLK_4_442_SplitCLK_4_441(net624_c1,net624);
INTERCONNECT SplitCLK_4_441_AND2T_31_n43(net625_c1,net625);
INTERCONNECT SplitCLK_4_441_DFFT_169__FPB_n496(net626_c1,net626);
INTERCONNECT SplitCLK_0_440_NOTT_12_n24(net627_c1,net627);
INTERCONNECT SplitCLK_0_440_DFFT_173__FPB_n500(net628_c1,net628);
INTERCONNECT SplitCLK_4_439_SplitCLK_4_437(net629_c1,net629);
INTERCONNECT SplitCLK_4_439_SplitCLK_4_438(net630_c1,net630);
INTERCONNECT SplitCLK_4_438_AND2T_17_n29(net631_c1,net631);
INTERCONNECT SplitCLK_4_438_AND2T_50_n62(net632_c1,net632);
INTERCONNECT SplitCLK_4_437_AND2T_134_n161(net633_c1,net633);
INTERCONNECT SplitCLK_4_437_AND2T_34_n46(net634_c1,net634);
INTERCONNECT SplitCLK_6_436_SplitCLK_6_405(net635_c1,net635);
INTERCONNECT SplitCLK_6_436_SplitCLK_2_435(net636_c1,net636);
INTERCONNECT SplitCLK_2_435_SplitCLK_6_420(net637_c1,net637);
INTERCONNECT SplitCLK_2_435_SplitCLK_4_434(net638_c1,net638);
INTERCONNECT SplitCLK_4_434_SplitCLK_6_427(net639_c1,net639);
INTERCONNECT SplitCLK_4_434_SplitCLK_2_433(net640_c1,net640);
INTERCONNECT SplitCLK_2_433_SplitCLK_6_430(net641_c1,net641);
INTERCONNECT SplitCLK_2_433_SplitCLK_4_432(net642_c1,net642);
INTERCONNECT SplitCLK_4_432_SplitCLK_4_500(net643_c1,net643);
INTERCONNECT SplitCLK_4_432_SplitCLK_4_431(net644_c1,net644);
INTERCONNECT SplitCLK_4_431_AND2T_56_n68(net645_c1,net645);
INTERCONNECT SplitCLK_4_431_AND2T_74_n86(net646_c1,net646);
INTERCONNECT SplitCLK_6_430_SplitCLK_4_428(net647_c1,net647);
INTERCONNECT SplitCLK_6_430_SplitCLK_4_429(net648_c1,net648);
INTERCONNECT SplitCLK_4_429_OR2T_76_n88(net649_c1,net649);
INTERCONNECT SplitCLK_4_429_OR2T_79_n91(net650_c1,net650);
INTERCONNECT SplitCLK_4_428_OR2T_66_n78(net651_c1,net651);
INTERCONNECT SplitCLK_4_428_OR2T_77_n89(net652_c1,net652);
INTERCONNECT SplitCLK_6_427_SplitCLK_4_423(net653_c1,net653);
INTERCONNECT SplitCLK_6_427_SplitCLK_4_426(net654_c1,net654);
INTERCONNECT SplitCLK_4_426_SplitCLK_4_424(net655_c1,net655);
INTERCONNECT SplitCLK_4_426_SplitCLK_4_425(net656_c1,net656);
INTERCONNECT SplitCLK_4_425_AND2T_51_n63(net657_c1,net657);
INTERCONNECT SplitCLK_4_425_OR2T_73_n85(net658_c1,net658);
INTERCONNECT SplitCLK_4_424_AND2T_25_n37(net659_c1,net659);
INTERCONNECT SplitCLK_4_424_OR2T_26_n38(net660_c1,net660);
INTERCONNECT SplitCLK_4_423_SplitCLK_0_421(net661_c1,net661);
INTERCONNECT SplitCLK_4_423_SplitCLK_4_422(net662_c1,net662);
INTERCONNECT SplitCLK_4_422_OR2T_59_n71(net663_c1,net663);
INTERCONNECT SplitCLK_4_422_OR2T_67_n79(net664_c1,net664);
INTERCONNECT SplitCLK_0_421_AND2T_60_n72(net665_c1,net665);
INTERCONNECT SplitCLK_0_421_DFFT_196__FPB_n523(net666_c1,net666);
INTERCONNECT SplitCLK_6_420_SplitCLK_6_412(net667_c1,net667);
INTERCONNECT SplitCLK_6_420_SplitCLK_2_419(net668_c1,net668);
INTERCONNECT SplitCLK_2_419_SplitCLK_2_415(net669_c1,net669);
INTERCONNECT SplitCLK_2_419_SplitCLK_4_418(net670_c1,net670);
INTERCONNECT SplitCLK_4_418_SplitCLK_4_416(net671_c1,net671);
INTERCONNECT SplitCLK_4_418_SplitCLK_4_417(net672_c1,net672);
INTERCONNECT SplitCLK_4_417_OR2T_58_n70(net673_c1,net673);
INTERCONNECT SplitCLK_4_417_DFFT_190__FPB_n517(net674_c1,net674);
INTERCONNECT SplitCLK_4_416_OR2T_68_n80(net675_c1,net675);
INTERCONNECT SplitCLK_4_416_DFFT_197__FPB_n524(net676_c1,net676);
INTERCONNECT SplitCLK_2_415_SplitCLK_4_413(net677_c1,net677);
INTERCONNECT SplitCLK_2_415_SplitCLK_4_414(net678_c1,net678);
INTERCONNECT SplitCLK_4_414_DFFT_143__FPB_n185(net679_c1,net679);
INTERCONNECT SplitCLK_4_414_DFFT_189__FPB_n516(net680_c1,net680);
INTERCONNECT SplitCLK_4_413_NOTT_49_n61(net681_c1,net681);
INTERCONNECT SplitCLK_4_413_DFFT_234__FPB_n561(net682_c1,net682);
INTERCONNECT SplitCLK_6_412_SplitCLK_0_408(net683_c1,net683);
INTERCONNECT SplitCLK_6_412_SplitCLK_4_411(net684_c1,net684);
INTERCONNECT SplitCLK_4_411_SplitCLK_4_409(net685_c1,net685);
INTERCONNECT SplitCLK_4_411_SplitCLK_4_410(net686_c1,net686);
INTERCONNECT SplitCLK_4_410_AND2T_114_n126(net687_c1,net687);
INTERCONNECT SplitCLK_4_410_AND2T_62_n74(net688_c1,net688);
INTERCONNECT SplitCLK_4_409_DFFT_207__FPB_n534(net689_c1,net689);
INTERCONNECT SplitCLK_4_409_DFFT_192__FPB_n519(net690_c1,net690);
INTERCONNECT SplitCLK_0_408_SplitCLK_4_406(net691_c1,net691);
INTERCONNECT SplitCLK_0_408_SplitCLK_0_407(net692_c1,net692);
INTERCONNECT SplitCLK_0_407_NOTT_138_n165(net693_c1,net693);
INTERCONNECT SplitCLK_0_407_DFFT_193__FPB_n520(net694_c1,net694);
INTERCONNECT SplitCLK_4_406_DFFT_204__FPB_n531(net695_c1,net695);
INTERCONNECT SplitCLK_4_406_DFFT_212__FPB_n539(net696_c1,net696);
INTERCONNECT SplitCLK_6_405_SplitCLK_6_389(net697_c1,net697);
INTERCONNECT SplitCLK_6_405_SplitCLK_4_404(net698_c1,net698);
INTERCONNECT SplitCLK_4_404_SplitCLK_0_396(net699_c1,net699);
INTERCONNECT SplitCLK_4_404_SplitCLK_2_403(net700_c1,net700);
INTERCONNECT SplitCLK_2_403_SplitCLK_2_399(net701_c1,net701);
INTERCONNECT SplitCLK_2_403_SplitCLK_2_402(net702_c1,net702);
INTERCONNECT SplitCLK_2_402_SplitCLK_4_400(net703_c1,net703);
INTERCONNECT SplitCLK_2_402_SplitCLK_4_401(net704_c1,net704);
INTERCONNECT SplitCLK_4_401_AND2T_85_n97(net705_c1,net705);
INTERCONNECT SplitCLK_4_401_OR2T_53_n65(net706_c1,net706);
INTERCONNECT SplitCLK_4_400_AND2T_75_n87(net707_c1,net707);
INTERCONNECT SplitCLK_4_400_OR2T_78_n90(net708_c1,net708);
INTERCONNECT SplitCLK_2_399_SplitCLK_4_397(net709_c1,net709);
INTERCONNECT SplitCLK_2_399_SplitCLK_4_398(net710_c1,net710);
INTERCONNECT SplitCLK_4_398_OR2T_55_n67(net711_c1,net711);
INTERCONNECT SplitCLK_4_398_DFFT_191__FPB_n518(net712_c1,net712);
INTERCONNECT SplitCLK_4_397_AND2T_61_n73(net713_c1,net713);
INTERCONNECT SplitCLK_4_397_OR2T_30_n42(net714_c1,net714);
INTERCONNECT SplitCLK_0_396_SplitCLK_6_392(net715_c1,net715);
INTERCONNECT SplitCLK_0_396_SplitCLK_4_395(net716_c1,net716);
INTERCONNECT SplitCLK_4_395_SplitCLK_4_393(net717_c1,net717);
INTERCONNECT SplitCLK_4_395_SplitCLK_4_394(net718_c1,net718);
INTERCONNECT SplitCLK_4_394_AND2T_28_n40(net719_c1,net719);
INTERCONNECT SplitCLK_4_394_NOTT_32_n44(net720_c1,net720);
INTERCONNECT SplitCLK_4_393_AND2T_84_n96(net721_c1,net721);
INTERCONNECT SplitCLK_4_393_DFFT_208__FPB_n535(net722_c1,net722);
INTERCONNECT SplitCLK_6_392_SplitCLK_4_390(net723_c1,net723);
INTERCONNECT SplitCLK_6_392_SplitCLK_4_391(net724_c1,net724);
INTERCONNECT SplitCLK_4_391_OR2T_108_n120(net725_c1,net725);
INTERCONNECT SplitCLK_4_391_DFFT_168__FPB_n495(net726_c1,net726);
INTERCONNECT SplitCLK_4_390_OR2T_109_n121(net727_c1,net727);
INTERCONNECT SplitCLK_4_390_DFFT_209__FPB_n536(net728_c1,net728);
INTERCONNECT SplitCLK_6_389_SplitCLK_6_381(net729_c1,net729);
INTERCONNECT SplitCLK_6_389_SplitCLK_6_388(net730_c1,net730);
INTERCONNECT SplitCLK_6_388_SplitCLK_6_384(net731_c1,net731);
INTERCONNECT SplitCLK_6_388_SplitCLK_4_387(net732_c1,net732);
INTERCONNECT SplitCLK_4_387_SplitCLK_4_385(net733_c1,net733);
INTERCONNECT SplitCLK_4_387_SplitCLK_4_386(net734_c1,net734);
INTERCONNECT SplitCLK_4_386_OR2T_69_n81(net735_c1,net735);
INTERCONNECT SplitCLK_4_386_AND2T_88_n100(net736_c1,net736);
INTERCONNECT SplitCLK_4_385_DFFT_210__FPB_n537(net737_c1,net737);
INTERCONNECT SplitCLK_4_385_OR2T_92_n104(net738_c1,net738);
INTERCONNECT SplitCLK_6_384_SplitCLK_4_382(net739_c1,net739);
INTERCONNECT SplitCLK_6_384_SplitCLK_4_383(net740_c1,net740);
INTERCONNECT SplitCLK_4_383_DFFT_213__FPB_n540(net741_c1,net741);
INTERCONNECT SplitCLK_4_383_DFFT_144__FPB_n186(net742_c1,net742);
INTERCONNECT SplitCLK_4_382_DFFT_214__FPB_n541(net743_c1,net743);
INTERCONNECT SplitCLK_4_382_DFFT_215__FPB_n542(net744_c1,net744);
INTERCONNECT SplitCLK_6_381_SplitCLK_0_377(net745_c1,net745);
INTERCONNECT SplitCLK_6_381_SplitCLK_4_380(net746_c1,net746);
INTERCONNECT SplitCLK_4_380_SplitCLK_4_378(net747_c1,net747);
INTERCONNECT SplitCLK_4_380_SplitCLK_4_379(net748_c1,net748);
INTERCONNECT SplitCLK_4_379_OR2T_115_n127(net749_c1,net749);
INTERCONNECT SplitCLK_4_379_DFFT_187__FPB_n514(net750_c1,net750);
INTERCONNECT SplitCLK_4_378_AND2T_112_n124(net751_c1,net751);
INTERCONNECT SplitCLK_4_378_DFFT_185__FPB_n512(net752_c1,net752);
INTERCONNECT SplitCLK_0_377_SplitCLK_4_375(net753_c1,net753);
INTERCONNECT SplitCLK_0_377_SplitCLK_0_376(net754_c1,net754);
INTERCONNECT SplitCLK_0_376_DFFT_242__FPB_n569(net755_c1,net755);
INTERCONNECT SplitCLK_0_376_DFFT_243__FPB_n570(net756_c1,net756);
INTERCONNECT SplitCLK_4_375_DFFT_205__FPB_n532(net757_c1,net757);
INTERCONNECT SplitCLK_4_375_DFFT_186__FPB_n513(net758_c1,net758);
INTERCONNECT SplitCLK_0_374_SplitCLK_6_312(net759_c1,net759);
INTERCONNECT SplitCLK_0_374_SplitCLK_4_373(net760_c1,net760);
INTERCONNECT SplitCLK_4_373_SplitCLK_0_342(net761_c1,net761);
INTERCONNECT SplitCLK_4_373_SplitCLK_4_372(net762_c1,net762);
INTERCONNECT SplitCLK_4_372_SplitCLK_6_357(net763_c1,net763);
INTERCONNECT SplitCLK_4_372_SplitCLK_4_371(net764_c1,net764);
INTERCONNECT SplitCLK_4_371_SplitCLK_0_364(net765_c1,net765);
INTERCONNECT SplitCLK_4_371_SplitCLK_6_370(net766_c1,net766);
INTERCONNECT SplitCLK_6_370_SplitCLK_6_367(net767_c1,net767);
INTERCONNECT SplitCLK_6_370_SplitCLK_6_369(net768_c1,net768);
INTERCONNECT SplitCLK_6_369_SplitCLK_2_499(net769_c1,net769);
INTERCONNECT SplitCLK_6_369_SplitCLK_4_368(net770_c1,net770);
INTERCONNECT SplitCLK_4_368_AND2T_137_n164(net771_c1,net771);
INTERCONNECT SplitCLK_4_368_DFFT_253__FPB_n580(net772_c1,net772);
INTERCONNECT SplitCLK_6_367_SplitCLK_4_365(net773_c1,net773);
INTERCONNECT SplitCLK_6_367_SplitCLK_4_366(net774_c1,net774);
INTERCONNECT SplitCLK_4_366_OR2T_18_n30(net775_c1,net775);
INTERCONNECT SplitCLK_4_366_OR2T_19_n31(net776_c1,net776);
INTERCONNECT SplitCLK_4_365_XOR2T_29_n41(net777_c1,net777);
INTERCONNECT SplitCLK_4_365_AND2T_37_n49(net778_c1,net778);
INTERCONNECT SplitCLK_0_364_SplitCLK_2_360(net779_c1,net779);
INTERCONNECT SplitCLK_0_364_SplitCLK_4_363(net780_c1,net780);
INTERCONNECT SplitCLK_4_363_SplitCLK_4_361(net781_c1,net781);
INTERCONNECT SplitCLK_4_363_SplitCLK_4_362(net782_c1,net782);
INTERCONNECT SplitCLK_4_362_DFFT_223__FPB_n550(net783_c1,net783);
INTERCONNECT SplitCLK_4_362_DFFT_155__FBL_n482(net784_c1,net784);
INTERCONNECT SplitCLK_4_361_DFFT_224__FPB_n551(net785_c1,net785);
INTERCONNECT SplitCLK_4_361_DFFT_225__FPB_n552(net786_c1,net786);
INTERCONNECT SplitCLK_2_360_SplitCLK_4_358(net787_c1,net787);
INTERCONNECT SplitCLK_2_360_SplitCLK_4_359(net788_c1,net788);
INTERCONNECT SplitCLK_4_359_AND2T_33_n45(net789_c1,net789);
INTERCONNECT SplitCLK_4_359_DFFT_227__FPB_n554(net790_c1,net790);
INTERCONNECT SplitCLK_4_358_AND2T_46_n58(net791_c1,net791);
INTERCONNECT SplitCLK_4_358_DFFT_170__FPB_n497(net792_c1,net792);
INTERCONNECT SplitCLK_6_357_SplitCLK_4_349(net793_c1,net793);
INTERCONNECT SplitCLK_6_357_SplitCLK_6_356(net794_c1,net794);
INTERCONNECT SplitCLK_6_356_SplitCLK_6_352(net795_c1,net795);
INTERCONNECT SplitCLK_6_356_SplitCLK_2_355(net796_c1,net796);
INTERCONNECT SplitCLK_2_355_SplitCLK_4_353(net797_c1,net797);
INTERCONNECT SplitCLK_2_355_SplitCLK_4_354(net798_c1,net798);
INTERCONNECT SplitCLK_4_354_OR2T_105_n117(net799_c1,net799);
INTERCONNECT SplitCLK_4_354_DFFT_174__FPB_n501(net800_c1,net800);
INTERCONNECT SplitCLK_4_353_DFFT_228__FPB_n555(net801_c1,net801);
INTERCONNECT SplitCLK_4_353_DFFT_176__FPB_n503(net802_c1,net802);
INTERCONNECT SplitCLK_6_352_SplitCLK_4_350(net803_c1,net803);
INTERCONNECT SplitCLK_6_352_SplitCLK_4_351(net804_c1,net804);
INTERCONNECT SplitCLK_4_351_NOTT_16_n28(net805_c1,net805);
INTERCONNECT SplitCLK_4_351_DFFT_175__FPB_n502(net806_c1,net806);
INTERCONNECT SplitCLK_4_350_DFFT_156__FBL_n483(net807_c1,net807);
INTERCONNECT SplitCLK_4_350_NOTT_142_n175(net808_c1,net808);
INTERCONNECT SplitCLK_4_349_SplitCLK_6_345(net809_c1,net809);
INTERCONNECT SplitCLK_4_349_SplitCLK_6_348(net810_c1,net810);
INTERCONNECT SplitCLK_6_348_SplitCLK_4_346(net811_c1,net811);
INTERCONNECT SplitCLK_6_348_SplitCLK_4_347(net812_c1,net812);
INTERCONNECT SplitCLK_4_347_AND2T_104_n116(net813_c1,net813);
INTERCONNECT SplitCLK_4_347_AND2T_48_n60(net814_c1,net814);
INTERCONNECT SplitCLK_4_346_AND2T_47_n59(net815_c1,net815);
INTERCONNECT SplitCLK_4_346_DFFT_177__FPB_n504(net816_c1,net816);
INTERCONNECT SplitCLK_6_345_SplitCLK_4_343(net817_c1,net817);
INTERCONNECT SplitCLK_6_345_SplitCLK_0_344(net818_c1,net818);
INTERCONNECT SplitCLK_0_344_AND2T_83_n95(net819_c1,net819);
INTERCONNECT SplitCLK_0_344_DFFT_149__FBL_n476(net820_c1,net820);
INTERCONNECT SplitCLK_4_343_OR2T_71_n83(net821_c1,net821);
INTERCONNECT SplitCLK_4_343_DFFT_145__FBL_n472(net822_c1,net822);
INTERCONNECT SplitCLK_0_342_SplitCLK_6_327(net823_c1,net823);
INTERCONNECT SplitCLK_0_342_SplitCLK_4_341(net824_c1,net824);
INTERCONNECT SplitCLK_4_341_SplitCLK_0_334(net825_c1,net825);
INTERCONNECT SplitCLK_4_341_SplitCLK_2_340(net826_c1,net826);
INTERCONNECT SplitCLK_2_340_SplitCLK_6_337(net827_c1,net827);
INTERCONNECT SplitCLK_2_340_SplitCLK_4_339(net828_c1,net828);
INTERCONNECT SplitCLK_4_339_SplitCLK_2_504(net829_c1,net829);
INTERCONNECT SplitCLK_4_339_SplitCLK_4_338(net830_c1,net830);
INTERCONNECT SplitCLK_4_338_DFFT_237__FPB_n564(net831_c1,net831);
INTERCONNECT SplitCLK_4_338_DFFT_238__FPB_n565(net832_c1,net832);
INTERCONNECT SplitCLK_6_337_SplitCLK_4_335(net833_c1,net833);
INTERCONNECT SplitCLK_6_337_SplitCLK_4_336(net834_c1,net834);
INTERCONNECT SplitCLK_4_336_AND2T_122_n134(net835_c1,net835);
INTERCONNECT SplitCLK_4_336_DFFT_241__FPB_n568(net836_c1,net836);
INTERCONNECT SplitCLK_4_335_AND2T_103_n115(net837_c1,net837);
INTERCONNECT SplitCLK_4_335_DFFT_163__FPB_n490(net838_c1,net838);
INTERCONNECT SplitCLK_0_334_SplitCLK_6_330(net839_c1,net839);
INTERCONNECT SplitCLK_0_334_SplitCLK_4_333(net840_c1,net840);
INTERCONNECT SplitCLK_4_333_SplitCLK_4_331(net841_c1,net841);
INTERCONNECT SplitCLK_4_333_SplitCLK_4_332(net842_c1,net842);
INTERCONNECT SplitCLK_4_332_DFFT_226__FPB_n553(net843_c1,net843);
INTERCONNECT SplitCLK_4_332_DFFT_239__FPB_n566(net844_c1,net844);
INTERCONNECT SplitCLK_4_331_AND2T_120_n132(net845_c1,net845);
INTERCONNECT SplitCLK_4_331_DFFT_240__FPB_n567(net846_c1,net846);
INTERCONNECT SplitCLK_6_330_SplitCLK_4_328(net847_c1,net847);
INTERCONNECT SplitCLK_6_330_SplitCLK_4_329(net848_c1,net848);
INTERCONNECT SplitCLK_4_329_AND2T_121_n133(net849_c1,net849);
INTERCONNECT SplitCLK_4_329_DFFT_221__FPB_n548(net850_c1,net850);
INTERCONNECT SplitCLK_4_328_AND2T_102_n114(net851_c1,net851);
INTERCONNECT SplitCLK_4_328_AND2T_97_n109(net852_c1,net852);
INTERCONNECT SplitCLK_6_327_SplitCLK_4_319(net853_c1,net853);
INTERCONNECT SplitCLK_6_327_SplitCLK_2_326(net854_c1,net854);
INTERCONNECT SplitCLK_2_326_SplitCLK_6_322(net855_c1,net855);
INTERCONNECT SplitCLK_2_326_SplitCLK_4_325(net856_c1,net856);
INTERCONNECT SplitCLK_4_325_SplitCLK_4_323(net857_c1,net857);
INTERCONNECT SplitCLK_4_325_SplitCLK_4_324(net858_c1,net858);
INTERCONNECT SplitCLK_4_324_OR2T_82_n94(net859_c1,net859);
INTERCONNECT SplitCLK_4_324_DFFT_178__FPB_n505(net860_c1,net860);
INTERCONNECT SplitCLK_4_323_AND2T_99_n111(net861_c1,net861);
INTERCONNECT SplitCLK_4_323_DFFT_203__FPB_n530(net862_c1,net862);
INTERCONNECT SplitCLK_6_322_SplitCLK_4_320(net863_c1,net863);
INTERCONNECT SplitCLK_6_322_SplitCLK_4_321(net864_c1,net864);
INTERCONNECT SplitCLK_4_321_DFFT_157__FBL_n484(net865_c1,net865);
INTERCONNECT SplitCLK_4_321_NOTT_141_n174(net866_c1,net866);
INTERCONNECT SplitCLK_4_320_OR2T_132_n144(net867_c1,net867);
INTERCONNECT SplitCLK_4_320_DFFT_251__FPB_n578(net868_c1,net868);
INTERCONNECT SplitCLK_4_319_SplitCLK_0_315(net869_c1,net869);
INTERCONNECT SplitCLK_4_319_SplitCLK_4_318(net870_c1,net870);
INTERCONNECT SplitCLK_4_318_SplitCLK_4_316(net871_c1,net871);
INTERCONNECT SplitCLK_4_318_SplitCLK_4_317(net872_c1,net872);
INTERCONNECT SplitCLK_4_317_AND2T_133_n145(net873_c1,net873);
INTERCONNECT SplitCLK_4_317_AND2T_98_n110(net874_c1,net874);
INTERCONNECT SplitCLK_4_316_DFFT_220__FPB_n547(net875_c1,net875);
INTERCONNECT SplitCLK_4_316_DFFT_219__FPB_n546(net876_c1,net876);
INTERCONNECT SplitCLK_0_315_SplitCLK_4_313(net877_c1,net877);
INTERCONNECT SplitCLK_0_315_SplitCLK_0_314(net878_c1,net878);
INTERCONNECT SplitCLK_0_314_OR2T_131_n143(net879_c1,net879);
INTERCONNECT SplitCLK_0_314_DFFT_151__FBL_n478(net880_c1,net880);
INTERCONNECT SplitCLK_4_313_DFFT_217__FPB_n544(net881_c1,net881);
INTERCONNECT SplitCLK_4_313_DFFT_218__FPB_n545(net882_c1,net882);
INTERCONNECT SplitCLK_6_312_SplitCLK_6_281(net883_c1,net883);
INTERCONNECT SplitCLK_6_312_SplitCLK_2_311(net884_c1,net884);
INTERCONNECT SplitCLK_2_311_SplitCLK_6_296(net885_c1,net885);
INTERCONNECT SplitCLK_2_311_SplitCLK_4_310(net886_c1,net886);
INTERCONNECT SplitCLK_4_310_SplitCLK_4_303(net887_c1,net887);
INTERCONNECT SplitCLK_4_310_SplitCLK_6_309(net888_c1,net888);
INTERCONNECT SplitCLK_6_309_SplitCLK_6_306(net889_c1,net889);
INTERCONNECT SplitCLK_6_309_SplitCLK_2_308(net890_c1,net890);
INTERCONNECT SplitCLK_2_308_SplitCLK_2_501(net891_c1,net891);
INTERCONNECT SplitCLK_2_308_SplitCLK_4_307(net892_c1,net892);
INTERCONNECT SplitCLK_4_307_DFFT_236__FPB_n563(net893_c1,net893);
INTERCONNECT SplitCLK_4_307_DFFT_247__FPB_n574(net894_c1,net894);
INTERCONNECT SplitCLK_6_306_SplitCLK_4_304(net895_c1,net895);
INTERCONNECT SplitCLK_6_306_SplitCLK_4_305(net896_c1,net896);
INTERCONNECT SplitCLK_4_305_OR2T_127_n139(net897_c1,net897);
INTERCONNECT SplitCLK_4_305_AND2T_89_n101(net898_c1,net898);
INTERCONNECT SplitCLK_4_304_AND2T_27_n39(net899_c1,net899);
INTERCONNECT SplitCLK_4_304_AND2T_64_n76(net900_c1,net900);
INTERCONNECT SplitCLK_4_303_SplitCLK_6_299(net901_c1,net901);
INTERCONNECT SplitCLK_4_303_SplitCLK_6_302(net902_c1,net902);
INTERCONNECT SplitCLK_6_302_SplitCLK_4_300(net903_c1,net903);
INTERCONNECT SplitCLK_6_302_SplitCLK_4_301(net904_c1,net904);
INTERCONNECT SplitCLK_4_301_AND2T_125_n137(net905_c1,net905);
INTERCONNECT SplitCLK_4_301_DFFT_166__FPB_n493(net906_c1,net906);
INTERCONNECT SplitCLK_4_300_OR2T_126_n138(net907_c1,net907);
INTERCONNECT SplitCLK_4_300_DFFT_150__FBL_n477(net908_c1,net908);
INTERCONNECT SplitCLK_6_299_SplitCLK_4_297(net909_c1,net909);
INTERCONNECT SplitCLK_6_299_SplitCLK_4_298(net910_c1,net910);
INTERCONNECT SplitCLK_4_298_DFFT_146__FBL_n473(net911_c1,net911);
INTERCONNECT SplitCLK_4_298_DFFT_195__FPB_n522(net912_c1,net912);
INTERCONNECT SplitCLK_4_297_OR2T_86_n98(net913_c1,net913);
INTERCONNECT SplitCLK_4_297_OR2T_139_n166(net914_c1,net914);
INTERCONNECT SplitCLK_6_296_SplitCLK_2_288(net915_c1,net915);
INTERCONNECT SplitCLK_6_296_SplitCLK_6_295(net916_c1,net916);
INTERCONNECT SplitCLK_6_295_SplitCLK_6_291(net917_c1,net917);
INTERCONNECT SplitCLK_6_295_SplitCLK_6_294(net918_c1,net918);
INTERCONNECT SplitCLK_6_294_SplitCLK_4_292(net919_c1,net919);
INTERCONNECT SplitCLK_6_294_SplitCLK_4_293(net920_c1,net920);
INTERCONNECT SplitCLK_4_293_AND2T_65_n77(net921_c1,net921);
INTERCONNECT SplitCLK_4_293_OR2T_91_n103(net922_c1,net922);
INTERCONNECT SplitCLK_4_292_OR2T_117_n129(net923_c1,net923);
INTERCONNECT SplitCLK_4_292_OR2T_90_n102(net924_c1,net924);
INTERCONNECT SplitCLK_6_291_SplitCLK_4_289(net925_c1,net925);
INTERCONNECT SplitCLK_6_291_SplitCLK_4_290(net926_c1,net926);
INTERCONNECT SplitCLK_4_290_OR2T_128_n140(net927_c1,net927);
INTERCONNECT SplitCLK_4_290_DFFT_232__FPB_n559(net928_c1,net928);
INTERCONNECT SplitCLK_4_289_DFFT_231__FPB_n558(net929_c1,net929);
INTERCONNECT SplitCLK_4_289_DFFT_181__FPB_n508(net930_c1,net930);
INTERCONNECT SplitCLK_2_288_SplitCLK_0_284(net931_c1,net931);
INTERCONNECT SplitCLK_2_288_SplitCLK_2_287(net932_c1,net932);
INTERCONNECT SplitCLK_2_287_SplitCLK_4_285(net933_c1,net933);
INTERCONNECT SplitCLK_2_287_SplitCLK_4_286(net934_c1,net934);
INTERCONNECT SplitCLK_4_286_OR2T_116_n128(net935_c1,net935);
INTERCONNECT SplitCLK_4_286_DFFT_235__FPB_n562(net936_c1,net936);
INTERCONNECT SplitCLK_4_285_AND2T_106_n118(net937_c1,net937);
INTERCONNECT SplitCLK_4_285_DFFT_183__FPB_n510(net938_c1,net938);
INTERCONNECT SplitCLK_0_284_SplitCLK_4_282(net939_c1,net939);
INTERCONNECT SplitCLK_0_284_SplitCLK_0_283(net940_c1,net940);
INTERCONNECT SplitCLK_0_283_DFFT_206__FPB_n533(net941_c1,net941);
INTERCONNECT SplitCLK_0_283_DFFT_182__FPB_n509(net942_c1,net942);
INTERCONNECT SplitCLK_4_282_AND2T_87_n99(net943_c1,net943);
INTERCONNECT SplitCLK_4_282_DFFT_184__FPB_n511(net944_c1,net944);
INTERCONNECT SplitCLK_6_281_SplitCLK_6_265(net945_c1,net945);
INTERCONNECT SplitCLK_6_281_SplitCLK_4_280(net946_c1,net946);
INTERCONNECT SplitCLK_4_280_SplitCLK_4_272(net947_c1,net947);
INTERCONNECT SplitCLK_4_280_SplitCLK_2_279(net948_c1,net948);
INTERCONNECT SplitCLK_2_279_SplitCLK_6_275(net949_c1,net949);
INTERCONNECT SplitCLK_2_279_SplitCLK_4_278(net950_c1,net950);
INTERCONNECT SplitCLK_4_278_SplitCLK_4_276(net951_c1,net951);
INTERCONNECT SplitCLK_4_278_SplitCLK_4_277(net952_c1,net952);
INTERCONNECT SplitCLK_4_277_OR2T_81_n93(net953_c1,net953);
INTERCONNECT SplitCLK_4_277_OR2T_100_n112(net954_c1,net954);
INTERCONNECT SplitCLK_4_276_OR2T_101_n113(net955_c1,net955);
INTERCONNECT SplitCLK_4_276_AND2T_96_n108(net956_c1,net956);
INTERCONNECT SplitCLK_6_275_SplitCLK_0_273(net957_c1,net957);
INTERCONNECT SplitCLK_6_275_SplitCLK_4_274(net958_c1,net958);
INTERCONNECT SplitCLK_4_274_AND2T_107_n119(net959_c1,net959);
INTERCONNECT SplitCLK_4_274_DFFT_230__FPB_n557(net960_c1,net960);
INTERCONNECT SplitCLK_0_273_OR2T_70_n82(net961_c1,net961);
INTERCONNECT SplitCLK_0_273_DFFT_229__FPB_n556(net962_c1,net962);
INTERCONNECT SplitCLK_4_272_SplitCLK_6_268(net963_c1,net963);
INTERCONNECT SplitCLK_4_272_SplitCLK_0_271(net964_c1,net964);
INTERCONNECT SplitCLK_0_271_SplitCLK_4_269(net965_c1,net965);
INTERCONNECT SplitCLK_0_271_SplitCLK_4_270(net966_c1,net966);
INTERCONNECT SplitCLK_4_270_DFFT_199__FPB_n526(net967_c1,net967);
INTERCONNECT SplitCLK_4_270_AND2T_94_n106(net968_c1,net968);
INTERCONNECT SplitCLK_4_269_DFFT_200__FPB_n527(net969_c1,net969);
INTERCONNECT SplitCLK_4_269_DFFT_222__FPB_n549(net970_c1,net970);
INTERCONNECT SplitCLK_6_268_SplitCLK_4_266(net971_c1,net971);
INTERCONNECT SplitCLK_6_268_SplitCLK_4_267(net972_c1,net972);
INTERCONNECT SplitCLK_4_267_OR2T_80_n92(net973_c1,net973);
INTERCONNECT SplitCLK_4_267_DFFT_202__FPB_n529(net974_c1,net974);
INTERCONNECT SplitCLK_4_266_OR2T_111_n123(net975_c1,net975);
INTERCONNECT SplitCLK_4_266_AND2T_95_n107(net976_c1,net976);
INTERCONNECT SplitCLK_6_265_SplitCLK_4_257(net977_c1,net977);
INTERCONNECT SplitCLK_6_265_SplitCLK_2_264(net978_c1,net978);
INTERCONNECT SplitCLK_2_264_SplitCLK_0_260(net979_c1,net979);
INTERCONNECT SplitCLK_2_264_SplitCLK_2_263(net980_c1,net980);
INTERCONNECT SplitCLK_2_263_SplitCLK_4_261(net981_c1,net981);
INTERCONNECT SplitCLK_2_263_SplitCLK_4_262(net982_c1,net982);
INTERCONNECT SplitCLK_4_262_DFFT_211__FPB_n538(net983_c1,net983);
INTERCONNECT SplitCLK_4_262_OR2T_93_n105(net984_c1,net984);
INTERCONNECT SplitCLK_4_261_AND2T_110_n122(net985_c1,net985);
INTERCONNECT SplitCLK_4_261_DFFT_216__FPB_n543(net986_c1,net986);
INTERCONNECT SplitCLK_0_260_SplitCLK_4_258(net987_c1,net987);
INTERCONNECT SplitCLK_0_260_SplitCLK_0_259(net988_c1,net988);
INTERCONNECT SplitCLK_0_259_AND2T_124_n136(net989_c1,net989);
INTERCONNECT SplitCLK_0_259_DFFT_245__FPB_n572(net990_c1,net990);
INTERCONNECT SplitCLK_4_258_DFFT_246__FPB_n573(net991_c1,net991);
INTERCONNECT SplitCLK_4_258_DFFT_248__FPB_n575(net992_c1,net992);
INTERCONNECT SplitCLK_4_257_SplitCLK_0_253(net993_c1,net993);
INTERCONNECT SplitCLK_4_257_SplitCLK_6_256(net994_c1,net994);
INTERCONNECT SplitCLK_6_256_SplitCLK_4_254(net995_c1,net995);
INTERCONNECT SplitCLK_6_256_SplitCLK_4_255(net996_c1,net996);
INTERCONNECT SplitCLK_4_255_AND2T_54_n66(net997_c1,net997);
INTERCONNECT SplitCLK_4_255_OR2T_129_n141(net998_c1,net998);
INTERCONNECT SplitCLK_4_254_OR2T_130_n142(net999_c1,net999);
INTERCONNECT SplitCLK_4_254_DFFT_198__FPB_n525(net1000_c1,net1000);
INTERCONNECT SplitCLK_0_253_SplitCLK_4_251(net1001_c1,net1001);
INTERCONNECT SplitCLK_0_253_SplitCLK_0_252(net1002_c1,net1002);
INTERCONNECT SplitCLK_0_252_AND2T_123_n135(net1003_c1,net1003);
INTERCONNECT SplitCLK_0_252_DFFT_244__FPB_n571(net1004_c1,net1004);
INTERCONNECT SplitCLK_4_251_DFFT_250__FPB_n577(net1005_c1,net1005);
INTERCONNECT SplitCLK_4_251_DFFT_249__FPB_n576(net1006_c1,net1006);
INTERCONNECT GCLK_Pad_SplitCLK_0_505(GCLK_Pad,net1007);
INTERCONNECT Split_HOLD_635_DFFT_162__FPB_n489(net1008_c1,net1008);

endmodule
